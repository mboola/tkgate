//: version "1.8.7"

module half_adder;    //: root_module
wire w6;    //: /sn:0 {0}(217,298)(217,314)(262,314)(262,242){1}
wire w7;    //: /sn:0 {0}(201,201)(201,217)(239,217){1}
wire w4;    //: /sn:0 {0}(164,173)(252,173)(252,196){1}
wire w5;    //: /sn:0 {0}(257,138)(271,138)(271,196){1}
//: enddecls

  led g4 (.I(w7));   //: @(201,194) /sn:0 /w:[ 0 ] /type:0
  led g3 (.I(w6));   //: @(217,291) /sn:0 /w:[ 0 ] /type:0
  //: switch g2 (w5) @(240,138) /sn:0 /w:[ 0 ] /st:0
  //: switch g1 (w4) @(147,173) /sn:0 /w:[ 0 ] /st:0
  HA g0 (.b(w5), .a(w4), .c(w7), .s(w6));   //: @(240, 197) /sz:(44, 44) /sn:0 /p:[ Ti0>1 Ti1>1 Lo0<1 Bo0<1 ]

endmodule

module HA(s, b, a, c);
//: interface  /sz:(44, 44) /bd:[ Ti0>b(31/44) Ti1>a(12/44) Lo0<c(20/44) Bo0<s(22/44) ]
input b;    //: /sn:0 /dp:1 {0}(94,103)(125,103)(125,129){1}
//: {2}(127,131)(183,131){3}
//: {4}(125,133)(125,166)(183,166){5}
output s;    //: /sn:0 /dp:1 {0}(204,129)(241,129){1}
input a;    //: /sn:0 /dp:1 {0}(183,161)(137,161)(137,128){1}
//: {2}(139,126)(183,126){3}
//: {4}(137,124)(137,87)(95,87){5}
output c;    //: /sn:0 /dp:1 {0}(204,164)(243,164){1}
//: enddecls

  //: output g4 (s) @(238,129) /sn:0 /w:[ 1 ]
  //: input g3 (b) @(92,103) /sn:0 /w:[ 0 ]
  //: input g2 (a) @(93,87) /sn:0 /w:[ 5 ]
  and g1 (.I0(a), .I1(b), .Z(c));   //: @(194,164) /sn:0 /delay:" 5" /w:[ 0 5 0 ]
  //: joint g6 (b) @(125, 131) /w:[ 2 1 -1 4 ]
  //: joint g7 (a) @(137, 126) /w:[ 2 4 -1 1 ]
  //: output g5 (c) @(240,164) /sn:0 /w:[ 1 ]
  xor g0 (.I0(a), .I1(b), .Z(s));   //: @(194,129) /sn:0 /delay:" 6" /w:[ 3 3 0 ]

endmodule
