//: version "1.8.7"

module CSA(c_in, b, a, c_out, s);
//: interface  /sz:(129, 81) /bd:[ Ti0>b[3:0](86/129) Ti1>a[3:0](31/129) Ri0>c_in(40/81) Lo0<c_out(38/81) Bo0<s[3:0](65/129) ]
input [3:0] b;    //: /sn:0 /dp:5 {0}(566,312)(566,116){1}
//: {2}(568,114)(728,114)(728,200){3}
//: {4}(564,114)(218,114){5}
output c_out;    //: /sn:0 /dp:1 {0}(410,399)(410,559)(827,559){1}
input c_in;    //: /sn:0 {0}(532,468)(313,468)(313,388){1}
//: {2}(315,386)(387,386){3}
//: {4}(313,384)(313,80)(214,80){5}
output [3:0] s;    //: /sn:0 /dp:1 {0}(555,481)(555,536)(826,536){1}
input [3:0] a;    //: /sn:0 {0}(523,312)(523,143){1}
//: {2}(525,141)(685,141)(685,200){3}
//: {4}(521,141)(220,141){5}
wire w7;    //: /sn:0 {0}(590,353)(652,353)(652,324)(642,324){1}
wire [3:0] w4;    //: /sn:0 {0}(707,281)(707,442)(565,442)(565,452){1}
wire w3;    //: /sn:0 {0}(660,242)(400,242)(400,370){1}
wire w8;    //: /sn:0 {0}(498,354)(420,354)(420,370){1}
wire w2;    //: /sn:0 {0}(752,241)(830,241)(830,211)(808,211){1}
wire [3:0] w9;    //: /sn:0 {0}(545,393)(545,452){1}
//: enddecls

  //: input g4 (c_in) @(212,80) /sn:0 /w:[ 5 ]
  //: joint g8 (b) @(566, 114) /w:[ 2 -1 4 1 ]
  //: input g3 (b) @(216,114) /sn:0 /w:[ 5 ]
  //: input g2 (a) @(218,141) /sn:0 /w:[ 5 ]
  CPA g1 (.a(a), .b(b), .c_in(w7), .c_out(w8), .s(w9));   //: @(499, 313) /sz:(90, 79) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>0 Lo0<0 Bo0<0 ]
  mux g10 (.I0(w3), .I1(w8), .S(c_in), .Z(c_out));   //: @(410,386) /sn:0 /w:[ 1 1 3 0 ] /ss:0 /do:0
  //: switch g6 (w7) @(625,324) /sn:0 /w:[ 1 ] /st:1
  //: joint g7 (a) @(523, 141) /w:[ 2 -1 4 1 ]
  mux g9 (.I0(w4), .I1(w9), .S(c_in), .Z(s));   //: @(555,468) /sn:0 /w:[ 1 1 0 0 ] /ss:0 /do:1
  //: output g12 (c_out) @(824,559) /sn:0 /w:[ 1 ]
  //: switch g5 (w2) @(791,211) /sn:0 /w:[ 1 ] /st:0
  //: joint g11 (c_in) @(313, 386) /w:[ 2 4 -1 1 ]
  CPA g0 (.a(a), .b(b), .c_in(w2), .c_out(w3), .s(w4));   //: @(661, 201) /sz:(90, 79) /sn:0 /p:[ Ti0>3 Ti1>3 Ri0>0 Lo0<0 Bo0<0 ]
  //: output g13 (s) @(823,536) /sn:0 /w:[ 1 ]

endmodule

module CPA(c_out, s, c_in, b, a);
//: interface  /sz:(90, 79) /bd:[ Ti0>a[3:0](24/90) Ti1>b[3:0](67/90) Ri0>c_in(40/79) Lo0<c_out(41/79) Bo0<s[3:0](46/90) ]
input [3:0] b;    //: /sn:0 {0}(467,173)(428,173){1}
//: {2}(427,173)(342,173){3}
//: {4}(341,173)(257,173){5}
//: {6}(256,173)(170,173){7}
//: {8}(169,173)(90,173){9}
output c_out;    //: /sn:0 {0}(556,374)(138,374)(138,269)(148,269){1}
input c_in;    //: /sn:0 {0}(91,156)(499,156)(499,269)(465,269){1}
output [3:0] s;    //: /sn:0 /dp:1 {0}(512,336)(556,336){1}
input [3:0] a;    //: /sn:0 {0}(90,191)(189,191){1}
//: {2}(190,191)(276,191){3}
//: {4}(277,191)(361,191){5}
//: {6}(362,191)(447,191){7}
//: {8}(448,191)(466,191){9}
wire w16;    //: /sn:0 {0}(170,249)(170,177){1}
wire w6;    //: /sn:0 {0}(342,249)(342,177){1}
wire w4;    //: /sn:0 {0}(436,291)(436,351)(506,351){1}
wire w3;    //: /sn:0 {0}(406,269)(379,269){1}
wire w0;    //: /sn:0 {0}(448,249)(448,195){1}
wire w19;    //: /sn:0 {0}(178,291)(178,321)(506,321){1}
wire w12;    //: /sn:0 {0}(294,269)(320,269){1}
wire w10;    //: /sn:0 {0}(277,249)(277,195){1}
wire w1;    //: /sn:0 {0}(428,249)(428,177){1}
wire w17;    //: /sn:0 {0}(207,269)(235,269){1}
wire w14;    //: /sn:0 {0}(265,291)(265,331)(506,331){1}
wire w11;    //: /sn:0 {0}(257,249)(257,177){1}
wire w15;    //: /sn:0 {0}(190,249)(190,195){1}
wire w5;    //: /sn:0 {0}(362,249)(362,195){1}
wire w9;    //: /sn:0 {0}(350,291)(350,341)(506,341){1}
//: enddecls

  FA g8 (.b(w16), .a(w15), .c_in(w17), .c_out(c_out), .s(w19));   //: @(149, 250) /sz:(57, 40) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>0 Lo0<1 Bo0<0 ]
  //: output g4 (c_out) @(553,374) /sn:0 /w:[ 0 ]
  tran g16(.Z(w11), .I(b[2]));   //: @(257,171) /sn:0 /R:1 /w:[ 1 6 5 ] /ss:1
  //: output g3 (s) @(553,336) /sn:0 /w:[ 1 ]
  tran g17(.Z(w16), .I(b[3]));   //: @(170,171) /sn:0 /R:1 /w:[ 1 8 7 ] /ss:1
  //: input g2 (c_in) @(89,156) /sn:0 /w:[ 0 ]
  //: input g1 (b) @(88,173) /sn:0 /w:[ 9 ]
  tran g10(.Z(w0), .I(a[0]));   //: @(448,189) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  FA g6 (.b(w6), .a(w5), .c_in(w3), .c_out(w12), .s(w9));   //: @(321, 250) /sz:(57, 40) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<1 Bo0<0 ]
  concat g9 (.I0(w4), .I1(w9), .I2(w14), .I3(w19), .Z(s));   //: @(511,336) /sn:0 /w:[ 1 1 1 1 0 ] /dr:0
  FA g7 (.b(w11), .a(w10), .c_in(w12), .c_out(w17), .s(w14));   //: @(236, 250) /sz:(57, 40) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>0 Lo0<1 Bo0<0 ]
  tran g12(.Z(w10), .I(a[2]));   //: @(277,189) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  tran g14(.Z(w1), .I(b[0]));   //: @(428,171) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:1
  tran g11(.Z(w5), .I(a[1]));   //: @(362,189) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  FA g5 (.b(w1), .a(w0), .c_in(c_in), .c_out(w3), .s(w4));   //: @(407, 250) /sz:(57, 40) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<0 Bo0<0 ]
  tran g15(.Z(w6), .I(b[1]));   //: @(342,171) /sn:0 /R:1 /w:[ 1 4 3 ] /ss:1
  //: input g0 (a) @(88,191) /sn:0 /w:[ 0 ]
  tran g13(.Z(w15), .I(a[3]));   //: @(190,189) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1

endmodule

module main;    //: root_module
wire [4:0] w6;    //: /sn:0 /dp:1 {0}(726,336)(726,424)(600,424){1}
wire [3:0] w4;    //: /sn:0 {0}(498,357)(498,429)(594,429){1}
wire [3:0] w0;    //: /sn:0 /dp:1 {0}(464,274)(464,193)(370,193)(370,107){1}
wire w3;    //: /sn:0 {0}(432,313)(397,313)(397,419)(594,419){1}
wire [3:0] w1;    //: /sn:0 /dp:1 {0}(519,274)(519,145)(460,145)(460,69){1}
wire w5;    //: /sn:0 {0}(569,108)(605,108)(605,315)(563,315){1}
//: enddecls

  concat g4 (.I0(w4), .I1(w3), .Z(w6));   //: @(599,424) /sn:0 /w:[ 1 1 1 ] /dr:0
  //: switch g3 (w5) @(552,108) /sn:0 /w:[ 0 ] /st:1
  //: dip g2 (w1) @(460,59) /sn:0 /w:[ 1 ] /st:15
  //: dip g1 (w0) @(370,97) /sn:0 /w:[ 1 ] /st:15
  led g6 (.I(w6));   //: @(726,329) /sn:0 /w:[ 0 ] /type:2
  CSA g0 (.b(w1), .a(w0), .c_in(w5), .c_out(w3), .s(w4));   //: @(433, 275) /sz:(129, 81) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<0 Bo0<0 ]

endmodule

module FA(c_out, s, c_in, b, a);
//: interface  /sz:(57, 40) /bd:[ Ti0>a(41/57) Ti1>b(21/57) Ri0>c_in(19/40) Lo0<c_out(19/40) Bo0<s(29/57) ]
input b;    //: /sn:0 {0}(156,62)(193,62)(193,98){1}
//: {2}(195,100)(233,100){3}
//: {4}(193,102)(193,162)(284,162){5}
output c_out;    //: /sn:0 /dp:1 {0}(366,145)(394,145){1}
input c_in;    //: /sn:0 /dp:1 {0}(156,46)(209,46)(209,116){1}
//: {2}(211,118)(327,118)(327,103)(344,103){3}
//: {4}(209,120)(209,144)(284,144){5}
output s;    //: /sn:0 /dp:1 {0}(365,101)(394,101){1}
input a;    //: /sn:0 {0}(156,78)(177,78)(177,93){1}
//: {2}(179,95)(233,95){3}
//: {4}(177,97)(177,167)(284,167){5}
wire w14;    //: /sn:0 {0}(305,165)(328,165)(328,147)(345,147){1}
wire w2;    //: /sn:0 {0}(254,98)(269,98){1}
//: {2}(273,98)(344,98){3}
//: {4}(271,100)(271,139)(284,139){5}
wire w11;    //: /sn:0 {0}(305,142)(345,142){1}
//: enddecls

  //: output g4 (c_out) @(391,145) /sn:0 /w:[ 1 ]
  and g8 (.I0(w2), .I1(c_in), .Z(w11));   //: @(295,142) /sn:0 /w:[ 5 5 0 ]
  //: output g3 (s) @(391,101) /sn:0 /w:[ 1 ]
  //: input g2 (c_in) @(154,46) /sn:0 /w:[ 0 ]
  //: input g1 (b) @(154,62) /sn:0 /w:[ 0 ]
  //: joint g10 (c_in) @(209, 118) /w:[ 2 1 -1 4 ]
  xor g6 (.I0(w2), .I1(c_in), .Z(s));   //: @(355,101) /sn:0 /w:[ 3 3 0 ]
  or g7 (.I0(w11), .I1(w14), .Z(c_out));   //: @(356,145) /sn:0 /w:[ 1 1 0 ]
  and g9 (.I0(b), .I1(a), .Z(w14));   //: @(295,165) /sn:0 /w:[ 5 5 0 ]
  //: joint g12 (b) @(193, 100) /w:[ 2 1 -1 4 ]
  //: joint g11 (w2) @(271, 98) /w:[ 2 -1 1 4 ]
  xor g5 (.I0(a), .I1(b), .Z(w2));   //: @(244,98) /sn:0 /w:[ 3 3 0 ]
  //: input g0 (a) @(154,78) /sn:0 /w:[ 0 ]
  //: joint g13 (a) @(177, 95) /w:[ 2 1 -1 4 ]

endmodule
