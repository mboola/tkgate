//: version "1.8.7"

module full_adder;    //: root_module
wire w4;    //: /sn:0 {0}(137,120)(137,137)(210,137){1}
wire w3;    //: /sn:0 {0}(178,186)(178,195)(240,195)(240,159){1}
wire w0;    //: /sn:0 {0}(179,22)(252,22)(252,117){1}
wire w1;    //: /sn:0 {0}(327,21)(337,21)(337,137)(269,137){1}
wire w5;    //: /sn:0 {0}(179,61)(232,61)(232,117){1}
//: enddecls

  led g4 (.I(w4));   //: @(137,113) /sn:0 /w:[ 0 ] /type:0
  //: switch g3 (w1) @(310,21) /sn:0 /w:[ 0 ] /st:0
  //: switch g2 (w0) @(162,22) /sn:0 /w:[ 0 ] /st:0
  //: switch g1 (w5) @(162,61) /sn:0 /w:[ 0 ] /st:0
  led g5 (.I(w3));   //: @(178,179) /sn:0 /w:[ 0 ] /type:0
  FA g0 (.a(w0), .b(w5), .c_in(w1), .c_out(w4), .s(w3));   //: @(211, 118) /sz:(57, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<1 Bo0<1 ]

endmodule

module FA(c_out, s, c_in, b, a);
//: interface  /sz:(57, 40) /bd:[ Ti0>b(21/57) Ti1>a(41/57) Ri0>c_in(19/40) Lo0<c_out(19/40) Bo0<s(29/57) ]
input b;    //: /sn:0 {0}(156,62)(193,62)(193,98){1}
//: {2}(195,100)(233,100){3}
//: {4}(193,102)(193,162)(284,162){5}
output c_out;    //: /sn:0 /dp:1 {0}(366,145)(394,145){1}
input c_in;    //: /sn:0 /dp:1 {0}(156,46)(209,46)(209,116){1}
//: {2}(211,118)(327,118)(327,103)(344,103){3}
//: {4}(209,120)(209,144)(284,144){5}
output s;    //: /sn:0 /dp:1 {0}(365,101)(394,101){1}
input a;    //: /sn:0 {0}(156,78)(177,78)(177,93){1}
//: {2}(179,95)(233,95){3}
//: {4}(177,97)(177,167)(284,167){5}
wire w14;    //: /sn:0 {0}(305,165)(328,165)(328,147)(345,147){1}
wire w11;    //: /sn:0 {0}(305,142)(345,142){1}
wire w2;    //: /sn:0 {0}(254,98)(269,98){1}
//: {2}(273,98)(344,98){3}
//: {4}(271,100)(271,139)(284,139){5}
//: enddecls

  and g8 (.I0(w2), .I1(c_in), .Z(w11));   //: @(295,142) /sn:0 /w:[ 5 5 0 ]
  //: output g4 (c_out) @(391,145) /sn:0 /w:[ 1 ]
  //: output g3 (s) @(391,101) /sn:0 /w:[ 1 ]
  //: input g2 (c_in) @(154,46) /sn:0 /w:[ 0 ]
  //: input g1 (b) @(154,62) /sn:0 /w:[ 0 ]
  //: joint g10 (c_in) @(209, 118) /w:[ 2 1 -1 4 ]
  xor g6 (.I0(w2), .I1(c_in), .Z(s));   //: @(355,101) /sn:0 /w:[ 3 3 0 ]
  and g9 (.I0(b), .I1(a), .Z(w14));   //: @(295,165) /sn:0 /w:[ 5 5 0 ]
  or g7 (.I0(w11), .I1(w14), .Z(c_out));   //: @(356,145) /sn:0 /w:[ 1 1 0 ]
  //: joint g12 (b) @(193, 100) /w:[ 2 1 -1 4 ]
  xor g5 (.I0(a), .I1(b), .Z(w2));   //: @(244,98) /sn:0 /w:[ 3 3 0 ]
  //: joint g11 (w2) @(271, 98) /w:[ 2 -1 1 4 ]
  //: input g0 (a) @(154,78) /sn:0 /w:[ 0 ]
  //: joint g13 (a) @(177, 95) /w:[ 2 1 -1 4 ]

endmodule
