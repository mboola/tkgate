//: version "1.8.7"

module CPA16(c_out, s, c_in, b, a);
//: interface  /sz:(97, 64) /bd:[ Ti0>b[15:0](67/97) Ti1>a[15:0](25/97) Ri0>c_in(29/64) Lo0<c_out(30/64) Bo0<s[15:0](50/97) ]
input [15:0] b;    //: /sn:0 {0}(620,123)(592,123){1}
//: {2}(591,123)(469,123){3}
//: {4}(468,123)(348,123){5}
//: {6}(347,123)(228,123){7}
//: {8}(227,123)(82,123){9}
output c_out;    //: /sn:0 {0}(681,413)(101,413)(101,262)(160,262){1}
input c_in;    //: /sn:0 {0}(80,92)(641,92)(641,260)(616,260){1}
output [15:0] s;    //: /sn:0 /dp:1 {0}(650,365)(681,365){1}
input [15:0] a;    //: /sn:0 {0}(82,155)(184,155){1}
//: {2}(185,155)(304,155){3}
//: {4}(305,155)(425,155){5}
//: {6}(426,155)(548,155){7}
//: {8}(549,155)(618,155){9}
wire [3:0] w6;    //: /sn:0 {0}(426,220)(426,159){1}
wire [3:0] w16;    //: /sn:0 {0}(644,360)(327,360)(327,301){1}
wire [3:0] w7;    //: /sn:0 {0}(348,220)(348,127){1}
wire [3:0] w4;    //: /sn:0 {0}(571,300)(571,380)(644,380){1}
wire [3:0] w0;    //: /sn:0 {0}(592,219)(592,127){1}
wire w3;    //: /sn:0 {0}(524,261)(493,261){1}
wire [3:0] w18;    //: /sn:0 {0}(644,350)(207,350)(207,301){1}
wire [3:0] w10;    //: /sn:0 {0}(305,220)(305,159){1}
wire [3:0] w1;    //: /sn:0 {0}(549,219)(549,159){1}
wire w8;    //: /sn:0 {0}(401,261)(372,261){1}
wire [3:0] w14;    //: /sn:0 {0}(185,220)(185,159){1}
wire [3:0] w11;    //: /sn:0 {0}(228,220)(228,127){1}
wire w15;    //: /sn:0 {0}(252,261)(280,261){1}
wire [3:0] w5;    //: /sn:0 {0}(469,220)(469,127){1}
wire [3:0] w9;    //: /sn:0 {0}(448,301)(448,370)(644,370){1}
//: enddecls

  //: output g4 (c_out) @(678,413) /sn:0 /w:[ 0 ]
  CPA g8 (.a(w14), .b(w11), .c_in(w15), .c_out(c_out), .s(w18));   //: @(161, 221) /sz:(90, 79) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>0 Lo0<1 Bo0<1 ]
  //: output g3 (s) @(678,365) /sn:0 /w:[ 1 ]
  tran g16(.Z(w6), .I(a[7:4]));   //: @(426,153) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  tran g17(.Z(w14), .I(a[15:12]));   //: @(185,153) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  //: input g2 (c_in) @(78,92) /sn:0 /w:[ 0 ]
  //: input g1 (b) @(80,123) /sn:0 /w:[ 9 ]
  tran g10(.Z(w5), .I(b[7:4]));   //: @(469,121) /sn:0 /R:1 /w:[ 1 4 3 ] /ss:1
  CPA g6 (.a(w6), .b(w5), .c_in(w3), .c_out(w8), .s(w9));   //: @(402, 221) /sz:(90, 79) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<0 Bo0<0 ]
  CPA g7 (.a(w10), .b(w7), .c_in(w8), .c_out(w15), .s(w16));   //: @(281, 221) /sz:(90, 79) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<1 Bo0<1 ]
  concat g9 (.I0(w4), .I1(w9), .I2(w16), .I3(w18), .Z(s));   //: @(649,365) /sn:0 /w:[ 1 1 0 0 0 ] /dr:0
  tran g12(.Z(w7), .I(b[11:8]));   //: @(348,121) /sn:0 /R:1 /w:[ 1 6 5 ] /ss:1
  CPA g5 (.a(w1), .b(w0), .c_in(c_in), .c_out(w3), .s(w4));   //: @(525, 220) /sz:(90, 79) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<0 Bo0<0 ]
  tran g11(.Z(w0), .I(b[3:0]));   //: @(592,121) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:1
  tran g14(.Z(w1), .I(a[3:0]));   //: @(549,153) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  //: input g0 (a) @(80,155) /sn:0 /w:[ 0 ]
  tran g15(.Z(w10), .I(a[11:8]));   //: @(305,153) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  tran g13(.Z(w11), .I(b[15:12]));   //: @(228,121) /sn:0 /R:1 /w:[ 1 8 7 ] /ss:1

endmodule

module CPA(c_out, s, c_in, b, a);
//: interface  /sz:(90, 79) /bd:[ Ti0>a[3:0](24/90) Ti1>b[3:0](67/90) Ri0>c_in(40/79) Lo0<c_out(41/79) Bo0<s[3:0](46/90) ]
input [3:0] b;    //: /sn:0 {0}(467,173)(428,173){1}
//: {2}(427,173)(342,173){3}
//: {4}(341,173)(257,173){5}
//: {6}(256,173)(170,173){7}
//: {8}(169,173)(90,173){9}
output c_out;    //: /sn:0 {0}(556,374)(138,374)(138,269)(148,269){1}
input c_in;    //: /sn:0 {0}(91,156)(499,156)(499,269)(465,269){1}
output [3:0] s;    //: /sn:0 /dp:1 {0}(512,336)(556,336){1}
input [3:0] a;    //: /sn:0 {0}(90,191)(189,191){1}
//: {2}(190,191)(276,191){3}
//: {4}(277,191)(361,191){5}
//: {6}(362,191)(447,191){7}
//: {8}(448,191)(466,191){9}
wire w16;    //: /sn:0 {0}(170,249)(170,177){1}
wire w6;    //: /sn:0 {0}(342,249)(342,177){1}
wire w4;    //: /sn:0 {0}(436,291)(436,351)(506,351){1}
wire w3;    //: /sn:0 {0}(406,269)(379,269){1}
wire w0;    //: /sn:0 {0}(448,249)(448,195){1}
wire w19;    //: /sn:0 {0}(178,291)(178,321)(506,321){1}
wire w12;    //: /sn:0 {0}(294,269)(320,269){1}
wire w10;    //: /sn:0 {0}(277,249)(277,195){1}
wire w1;    //: /sn:0 {0}(428,249)(428,177){1}
wire w17;    //: /sn:0 {0}(207,269)(235,269){1}
wire w14;    //: /sn:0 {0}(265,291)(265,331)(506,331){1}
wire w11;    //: /sn:0 {0}(257,249)(257,177){1}
wire w15;    //: /sn:0 {0}(190,249)(190,195){1}
wire w5;    //: /sn:0 {0}(362,249)(362,195){1}
wire w9;    //: /sn:0 {0}(350,291)(350,341)(506,341){1}
//: enddecls

  FA g8 (.b(w16), .a(w15), .c_in(w17), .c_out(c_out), .s(w19));   //: @(149, 250) /sz:(57, 40) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>0 Lo0<1 Bo0<0 ]
  //: output g4 (c_out) @(553,374) /sn:0 /w:[ 0 ]
  tran g16(.Z(w11), .I(b[2]));   //: @(257,171) /sn:0 /R:1 /w:[ 1 6 5 ] /ss:1
  //: output g3 (s) @(553,336) /sn:0 /w:[ 1 ]
  tran g17(.Z(w16), .I(b[3]));   //: @(170,171) /sn:0 /R:1 /w:[ 1 8 7 ] /ss:1
  //: input g2 (c_in) @(89,156) /sn:0 /w:[ 0 ]
  //: input g1 (b) @(88,173) /sn:0 /w:[ 9 ]
  tran g10(.Z(w0), .I(a[0]));   //: @(448,189) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  FA g6 (.b(w6), .a(w5), .c_in(w3), .c_out(w12), .s(w9));   //: @(321, 250) /sz:(57, 40) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<1 Bo0<0 ]
  concat g9 (.I0(w4), .I1(w9), .I2(w14), .I3(w19), .Z(s));   //: @(511,336) /sn:0 /w:[ 1 1 1 1 0 ] /dr:0
  FA g7 (.b(w11), .a(w10), .c_in(w12), .c_out(w17), .s(w14));   //: @(236, 250) /sz:(57, 40) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>0 Lo0<1 Bo0<0 ]
  tran g12(.Z(w10), .I(a[2]));   //: @(277,189) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  tran g14(.Z(w1), .I(b[0]));   //: @(428,171) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:1
  tran g11(.Z(w5), .I(a[1]));   //: @(362,189) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  FA g5 (.b(w1), .a(w0), .c_in(c_in), .c_out(w3), .s(w4));   //: @(407, 250) /sz:(57, 40) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<0 Bo0<0 ]
  tran g15(.Z(w6), .I(b[1]));   //: @(342,171) /sn:0 /R:1 /w:[ 1 4 3 ] /ss:1
  //: input g0 (a) @(88,191) /sn:0 /w:[ 0 ]
  tran g13(.Z(w15), .I(a[3]));   //: @(190,189) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1

endmodule

module main;    //: root_module
wire [15:0] w6;    //: /sn:0 {0}(246,108)(246,177)(293,177)(293,275){1}
wire w4;    //: /sn:0 {0}(225,303)(187,303)(187,379)(390,379){1}
wire w0;    //: /sn:0 {0}(314,135)(342,135)(342,302)(324,302){1}
wire [15:0] w1;    //: /sn:0 {0}(390,389)(276,389)(276,336){1}
wire [16:0] w2;    //: /sn:0 /dp:1 {0}(453,242)(453,384)(396,384){1}
wire [15:0] w5;    //: /sn:0 {0}(187,165)(187,216)(251,216)(251,275){1}
//: enddecls

  concat g4 (.I0(w1), .I1(w4), .Z(w2));   //: @(395,384) /sn:0 /w:[ 0 1 1 ] /dr:0
  //: switch g3 (w0) @(297,135) /sn:0 /w:[ 0 ] /st:1
  //: dip g2 (w6) @(246,98) /sn:0 /w:[ 0 ] /st:7
  //: dip g1 (w5) @(187,155) /sn:0 /w:[ 0 ] /st:7
  led g5 (.I(w2));   //: @(453,235) /sn:0 /w:[ 0 ] /type:1
  CPA16 g0 (.b(w6), .a(w5), .c_in(w0), .c_out(w4), .s(w1));   //: @(226, 276) /sz:(97, 59) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<1 ]

endmodule

module FA(c_out, s, c_in, b, a);
//: interface  /sz:(57, 40) /bd:[ Ti0>a(41/57) Ti1>b(21/57) Ri0>c_in(19/40) Lo0<c_out(19/40) Bo0<s(29/57) ]
input b;    //: /sn:0 {0}(49,62)(111,62){1}
output c_out;    //: /sn:0 /dp:1 {0}(366,145)(394,145){1}
input c_in;    //: /sn:0 /dp:1 {0}(156,46)(209,46)(209,116){1}
//: {2}(211,118)(327,118)(327,103)(344,103){3}
//: {4}(209,120)(209,144)(284,144){5}
output s;    //: /sn:0 /dp:1 {0}(365,101)(394,101){1}
input a;    //: /sn:0 {0}(156,78)(177,78)(177,93){1}
//: {2}(179,95)(233,95){3}
//: {4}(177,97)(177,167)(284,167){5}
wire w4;    //: /sn:0 {0}(132,65)(193,65)(193,98){1}
//: {2}(195,100)(233,100){3}
//: {4}(193,102)(193,162)(284,162){5}
wire w0;    //: /sn:0 {0}(79,121)(101,121)(101,67)(111,67){1}
wire w14;    //: /sn:0 {0}(305,165)(328,165)(328,147)(345,147){1}
wire w2;    //: /sn:0 {0}(254,98)(269,98){1}
//: {2}(273,98)(344,98){3}
//: {4}(271,100)(271,139)(284,139){5}
wire w11;    //: /sn:0 {0}(305,142)(345,142){1}
//: enddecls

  //: output g4 (c_out) @(391,145) /sn:0 /w:[ 1 ]
  and g8 (.I0(w2), .I1(c_in), .Z(w11));   //: @(295,142) /sn:0 /w:[ 5 5 0 ]
  //: output g3 (s) @(391,101) /sn:0 /w:[ 1 ]
  //: input g2 (c_in) @(154,46) /sn:0 /w:[ 0 ]
  //: input g1 (b) @(47,62) /sn:0 /w:[ 0 ]
  //: joint g10 (c_in) @(209, 118) /w:[ 2 1 -1 4 ]
  xor g6 (.I0(w2), .I1(c_in), .Z(s));   //: @(355,101) /sn:0 /w:[ 3 3 0 ]
  or g7 (.I0(w11), .I1(w14), .Z(c_out));   //: @(356,145) /sn:0 /w:[ 1 1 0 ]
  and g9 (.I0(w4), .I1(a), .Z(w14));   //: @(295,165) /sn:0 /w:[ 5 5 0 ]
  xor g12 (.I0(b), .I1(w0), .Z(w4));   //: @(122,65) /sn:0 /w:[ 1 1 0 ]
  //: joint g14 (w4) @(193, 100) /w:[ 2 1 -1 4 ]
  //: joint g11 (w2) @(271, 98) /w:[ 2 -1 1 4 ]
  xor g5 (.I0(a), .I1(w4), .Z(w2));   //: @(244,98) /sn:0 /w:[ 3 3 0 ]
  //: switch g15 (w0) @(62,121) /sn:0 /w:[ 0 ] /st:1
  //: input g0 (a) @(154,78) /sn:0 /w:[ 0 ]
  //: joint g13 (a) @(177, 95) /w:[ 2 1 -1 4 ]

endmodule
