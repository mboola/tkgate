//: version "1.8.7"

module half_adder;    //: root_module
wire w6;    //: /sn:0 {0}(217,298)(217,314)(262,314)(262,242){1}
wire w7;    //: /sn:0 {0}(201,201)(201,217)(239,217){1}
wire w4;    //: /sn:0 {0}(164,173)(252,173)(252,196){1}
wire w5;    //: /sn:0 {0}(257,138)(271,138)(271,196){1}
//: enddecls

  led g4 (.I(w7));   //: @(201,194) /sn:0 /w:[ 0 ] /type:0
  led g3 (.I(w6));   //: @(217,291) /sn:0 /w:[ 0 ] /type:0
  //: switch g2 (w5) @(240,138) /sn:0 /w:[ 0 ] /st:0
  //: switch g1 (w4) @(147,173) /sn:0 /w:[ 0 ] /st:0
  HA g0 (.b(w5), .a(w4), .c(w7), .s(w6));   //: @(240, 197) /sz:(44, 44) /sn:0 /p:[ Ti0>1 Ti1>1 Lo0<1 Bo0<1 ]

endmodule

module HA(s, b, a, c);
//: interface  /sz:(44, 44) /bd:[ Ti0>a(11/40) Ti1>b(29/40) Lo0<c(19/40) Bo0<s(20/40) ]
input b;    //: /sn:0 /dp:1 {0}(180,145)(134,145){1}
//: {2}(132,143)(132,102)(180,102){3}
//: {4}(130,145)(91,145){5}
output s;    //: /sn:0 /dp:1 {0}(201,100)(238,100){1}
input a;    //: /sn:0 /dp:1 {0}(180,140)(151,140)(151,99){1}
//: {2}(153,97)(180,97){3}
//: {4}(149,97)(90,97){5}
output c;    //: /sn:0 /dp:1 {0}(201,143)(240,143){1}
//: enddecls

  //: output g4 (s) @(235,100) /sn:0 /w:[ 1 ]
  //: input g3 (b) @(89,145) /sn:0 /w:[ 5 ]
  //: input g2 (a) @(88,97) /sn:0 /w:[ 5 ]
  and g1 (.I0(a), .I1(b), .Z(c));   //: @(191,143) /sn:0 /delay:" 5" /w:[ 0 0 0 ]
  //: joint g6 (b) @(132, 145) /w:[ 1 2 4 -1 ]
  //: joint g7 (a) @(151, 97) /w:[ 2 -1 4 1 ]
  //: output g5 (c) @(237,143) /sn:0 /w:[ 1 ]
  xor g0 (.I0(a), .I1(b), .Z(s));   //: @(191,100) /sn:0 /delay:" 6" /w:[ 3 3 0 ]

endmodule
