//: version "1.8.7"

module PFA(p, c, b, s, g, a);
//: interface  /sz:(52, 50) /bd:[ Ti0>b(36/52) Ti1>a(14/52) Ri0>c(26/50) Bo0<p(9/52) Bo1<g(25/52) Bo2<s(41/52) ]
output p;    //: /sn:0 {0}(506,190)(454,190){1}
input b;    //: /sn:0 {0}(265,98)(265,147){1}
//: {2}(267,149)(341,149){3}
//: {4}(265,151)(265,190){5}
//: {6}(267,192)(433,192){7}
//: {8}(265,194)(265,222)(432,222){9}
output s;    //: /sn:0 /dp:1 {0}(453,159)(506,159){1}
input a;    //: /sn:0 {0}(291,98)(291,142){1}
//: {2}(293,144)(341,144){3}
//: {4}(291,146)(291,185){5}
//: {6}(293,187)(433,187){7}
//: {8}(291,189)(291,217)(432,217){9}
input c;    //: /sn:0 {0}(242,98)(242,161)(432,161){1}
output g;    //: /sn:0 {0}(506,220)(453,220){1}
wire w2;    //: /sn:0 {0}(362,147)(393,147)(393,156)(432,156){1}
//: enddecls

  xor g4 (.I0(w2), .I1(c), .Z(s));   //: @(443,159) /sn:0 /delay:" 6" /w:[ 1 1 0 ]
  //: output g8 (p) @(503,190) /sn:0 /w:[ 0 ]
  xor g3 (.I0(a), .I1(b), .Z(w2));   //: @(352,147) /sn:0 /delay:" 6" /w:[ 3 3 0 ]
  //: input g2 (c) @(242,96) /sn:0 /R:3 /w:[ 0 ]
  //: input g1 (b) @(265,96) /sn:0 /R:3 /w:[ 0 ]
  //: joint g10 (a) @(291, 144) /w:[ 2 1 -1 4 ]
  and g6 (.I0(a), .I1(b), .Z(g));   //: @(443,220) /sn:0 /delay:" 5" /w:[ 9 9 1 ]
  //: output g7 (s) @(503,159) /sn:0 /w:[ 1 ]
  //: output g9 (g) @(503,220) /sn:0 /w:[ 0 ]
  //: joint g12 (a) @(291, 187) /w:[ 6 5 -1 8 ]
  or g5 (.I0(a), .I1(b), .Z(p));   //: @(444,190) /sn:0 /delay:" 5" /w:[ 7 7 1 ]
  //: joint g11 (b) @(265, 192) /w:[ 6 5 -1 8 ]
  //: input g0 (a) @(291,96) /sn:0 /R:3 /w:[ 0 ]
  //: joint g13 (b) @(265, 149) /w:[ 2 1 -1 4 ]

endmodule

module CarryLookaheadLogic(p3, g3, g2, g1, c3, c2, g0, p1, p2, c4, c1, p0, c0);
//: interface  /sz:(266, 40) /bd:[ Ti0>g0(239/266) Ti1>p0(223/266) Ti2>g1(168/266) Ti3>p1(152/266) Ti4>g2(96/266) Ti5>p2(80/266) Ti6>g3(25/266) Ti7>p3(9/266) Ri0>c0(20/40) To0<c1(204/266) To1<c2(133/266) To2<c3(62/266) Lo0<c4(19/41) ]
input g3;    //: /sn:0 {0}(183,69)(183,579)(278,579)(278,511)(306,511){1}
input g2;    //: /sn:0 {0}(286,338)(266,338)(266,359)(163,359){1}
//: {2}(161,357)(161,69){3}
//: {4}(161,361)(161,535)(219,535){5}
input c0;    //: /sn:0 /dp:11 {0}(221,278)(9,278){1}
//: {2}(7,276)(7,181){3}
//: {4}(9,179)(220,179){5}
//: {6}(7,177)(7,118){7}
//: {8}(9,116)(220,116){9}
//: {10}(7,114)(7,69){11}
//: {12}(7,280)(7,403)(221,403){13}
input g1;    //: /sn:0 {0}(221,348)(142,348){1}
//: {2}(140,346)(140,240){3}
//: {4}(142,238)(253,238)(253,224)(287,224){5}
//: {6}(140,236)(140,69){7}
//: {8}(140,350)(140,506)(219,506){9}
output c4;    //: /sn:0 {0}(362,501)(327,501){1}
output c1;    //: /sn:0 {0}(359,128)(308,128){1}
input p3;    //: /sn:0 {0}(220,464)(90,464){1}
//: {2}(88,462)(88,425){3}
//: {4}(90,423)(221,423){5}
//: {6}(88,421)(88,69){7}
//: {8}(88,466)(88,499){9}
//: {10}(90,501)(219,501){11}
//: {12}(88,503)(88,530)(219,530){13}
input p2;    //: /sn:0 {0}(221,418)(71,418){1}
//: {2}(69,416)(69,345){3}
//: {4}(71,343)(221,343){5}
//: {6}(69,341)(69,321){7}
//: {8}(71,319)(221,319){9}
//: {10}(69,317)(69,295){11}
//: {12}(71,293)(221,293){13}
//: {14}(69,291)(69,69){15}
//: {16}(69,420)(69,457){17}
//: {18}(71,459)(220,459){19}
//: {20}(69,461)(69,496)(219,496){21}
output c3;    //: /sn:0 {0}(361,330)(307,330){1}
input p1;    //: /sn:0 {0}(221,413)(52,413){1}
//: {2}(50,411)(50,316){3}
//: {4}(52,314)(221,314){5}
//: {6}(50,312)(50,290){7}
//: {8}(52,288)(221,288){9}
//: {10}(50,286)(50,218){11}
//: {12}(52,216)(220,216){13}
//: {14}(50,214)(50,191){15}
//: {16}(52,189)(220,189){17}
//: {18}(50,187)(50,69){19}
//: {20}(50,415)(50,454)(220,454){21}
input p0;    //: /sn:0 /dp:7 {0}(220,184)(34,184){1}
//: {2}(32,182)(32,123){3}
//: {4}(34,121)(220,121){5}
//: {6}(32,119)(32,69){7}
//: {8}(32,186)(32,281){9}
//: {10}(34,283)(221,283){11}
//: {12}(32,285)(32,408)(221,408){13}
output c2;    //: /sn:0 {0}(359,219)(308,219){1}
input g0;    //: /sn:0 {0}(221,324)(122,324){1}
//: {2}(120,322)(120,223){3}
//: {4}(122,221)(220,221){5}
//: {6}(120,219)(120,132){7}
//: {8}(122,130)(287,130){9}
//: {10}(120,128)(120,69){11}
//: {12}(120,326)(120,469)(220,469){13}
wire w16;    //: /sn:0 {0}(306,506)(261,506)(261,533)(240,533){1}
wire w4;    //: /sn:0 /dp:1 {0}(286,328)(256,328)(256,319)(242,319){1}
wire w0;    //: /sn:0 /dp:1 {0}(287,214)(253,214)(253,184)(241,184){1}
wire w3;    //: /sn:0 /dp:1 {0}(241,119)(251,119)(251,125)(287,125){1}
wire w12;    //: /sn:0 {0}(240,501)(306,501){1}
wire w1;    //: /sn:0 /dp:1 {0}(287,219)(241,219){1}
wire w8;    //: /sn:0 /dp:1 {0}(306,496)(259,496)(259,461)(241,461){1}
wire w2;    //: /sn:0 /dp:1 {0}(286,323)(266,323)(266,285)(242,285){1}
wire w5;    //: /sn:0 /dp:1 {0}(306,491)(276,491)(276,413)(242,413){1}
wire w9;    //: /sn:0 {0}(242,346)(256,346)(256,333)(286,333){1}
//: enddecls

  //: joint g44 (p2) @(69, 418) /w:[ 1 2 -1 16 ]
  //: input g8 (p3) @(88,67) /sn:0 /R:3 /w:[ 7 ]
  //: input g4 (g3) @(183,67) /sn:0 /R:3 /w:[ 0 ]
  //: joint g16 (c0) @(7, 179) /w:[ 4 6 -1 3 ]
  //: input g3 (g2) @(161,67) /sn:0 /R:3 /w:[ 3 ]
  //: joint g17 (p0) @(32, 184) /w:[ 1 2 -1 8 ]
  //: joint g26 (c0) @(7, 278) /w:[ 1 2 -1 12 ]
  //: input g2 (g1) @(140,67) /sn:0 /R:3 /w:[ 7 ]
  and g30 (.I0(p1), .I1(p2), .I2(g0), .Z(w4));   //: @(232,319) /sn:0 /delay:" 5" /w:[ 5 9 0 1 ]
  //: joint g23 (g1) @(140, 238) /w:[ 4 6 -1 3 ]
  //: output g39 (c3) @(358,330) /sn:0 /w:[ 0 ]
  //: output g24 (c2) @(356,219) /sn:0 /w:[ 0 ]
  //: input g1 (g0) @(120,67) /sn:0 /R:3 /w:[ 11 ]
  //: joint g29 (p2) @(69, 293) /w:[ 12 14 -1 11 ]
  and g51 (.I0(p2), .I1(p3), .I2(g1), .Z(w12));   //: @(230,501) /sn:0 /w:[ 21 11 9 0 ]
  //: joint g18 (p1) @(50, 189) /w:[ 16 18 -1 15 ]
  and g25 (.I0(c0), .I1(p0), .I2(p1), .I3(p2), .Z(w2));   //: @(232,285) /sn:0 /delay:" 5" /w:[ 0 11 9 13 1 ]
  or g10 (.I0(w3), .I1(g0), .Z(c1));   //: @(298,128) /sn:0 /delay:" 5" /w:[ 1 9 1 ]
  //: joint g49 (p3) @(88, 464) /w:[ 1 2 -1 8 ]
  //: input g6 (p1) @(50,67) /sn:0 /R:3 /w:[ 19 ]
  or g58 (.I0(w5), .I1(w8), .I2(w12), .I3(w16), .I4(g3), .Z(c4));   //: @(317,501) /sn:0 /w:[ 0 0 1 0 1 1 ]
  //: joint g35 (p2) @(69, 343) /w:[ 4 6 -1 3 ]
  and g9 (.I0(c0), .I1(p0), .Z(w3));   //: @(231,119) /sn:0 /delay:" 5" /w:[ 9 5 0 ]
  //: input g7 (p2) @(69,67) /sn:0 /R:3 /w:[ 15 ]
  //: joint g31 (p1) @(50, 314) /w:[ 4 6 -1 3 ]
  or g22 (.I0(w0), .I1(w1), .I2(g1), .Z(c2));   //: @(298,219) /sn:0 /delay:" 5" /w:[ 0 0 5 1 ]
  //: output g41 (c4) @(359,501) /sn:0 /w:[ 0 ]
  //: joint g45 (p3) @(88, 423) /w:[ 4 6 -1 3 ]
  //: joint g36 (g1) @(140, 348) /w:[ 1 2 -1 8 ]
  //: joint g33 (g0) @(120, 324) /w:[ 1 2 -1 12 ]
  and g40 (.I0(c0), .I1(p0), .I2(p1), .I3(p2), .I4(p3), .Z(w5));   //: @(232,413) /sn:0 /w:[ 13 13 0 0 5 1 ]
  //: joint g12 (p0) @(32, 121) /w:[ 4 6 -1 3 ]
  and g46 (.I0(p1), .I1(p2), .I2(p3), .I3(g0), .Z(w8));   //: @(231,461) /sn:0 /w:[ 21 19 0 13 1 ]
  and g34 (.I0(p2), .I1(g1), .Z(w9));   //: @(232,346) /sn:0 /delay:" 5" /w:[ 5 0 0 ]
  //: joint g28 (p1) @(50, 288) /w:[ 8 10 -1 7 ]
  //: joint g11 (c0) @(7, 116) /w:[ 8 10 -1 7 ]
  //: output g14 (c1) @(356,128) /sn:0 /w:[ 0 ]
  //: input g5 (p0) @(32,67) /sn:0 /R:3 /w:[ 7 ]
  //: joint g21 (g0) @(120, 221) /w:[ 4 6 -1 3 ]
  and g19 (.I0(p1), .I1(g0), .Z(w1));   //: @(231,219) /sn:0 /delay:" 5" /w:[ 13 5 1 ]
  //: joint g32 (p2) @(69, 319) /w:[ 8 10 -1 7 ]
  //: joint g20 (p1) @(50, 216) /w:[ 12 14 -1 11 ]
  //: joint g43 (p1) @(50, 413) /w:[ 1 2 -1 20 ]
  //: joint g38 (g2) @(161, 359) /w:[ 1 2 -1 4 ]
  and g15 (.I0(c0), .I1(p0), .I2(p1), .Z(w0));   //: @(231,184) /sn:0 /delay:" 5" /w:[ 5 0 17 1 ]
  //: input g0 (c0) @(7,67) /sn:0 /R:3 /w:[ 11 ]
  //: joint g48 (p2) @(69, 459) /w:[ 18 17 -1 20 ]
  //: joint g27 (p0) @(32, 283) /w:[ 10 9 -1 12 ]
  or g37 (.I0(w2), .I1(w4), .I2(w9), .I3(g2), .Z(c3));   //: @(297,330) /sn:0 /delay:" 5" /w:[ 0 0 1 0 1 ]
  and g55 (.I0(p3), .I1(g2), .Z(w16));   //: @(230,533) /sn:0 /w:[ 13 5 1 ]
  //: joint g53 (p3) @(88, 501) /w:[ 10 9 -1 12 ]
  //: joint g13 (g0) @(120, 130) /w:[ 8 10 -1 7 ]

endmodule

module main;    //: root_module
wire [3:0] w6;    //: /sn:0 {0}(484,156)(484,232)(450,232)(450,280){1}
wire w4;    //: /sn:0 {0}(406,310)(362,310){1}
wire [4:0] w0;    //: /sn:0 /dp:1 {0}(315,236)(315,305)(356,305){1}
wire [3:0] w3;    //: /sn:0 {0}(438,339)(438,358)(387,358)(387,300)(362,300){1}
wire w1;    //: /sn:0 {0}(514,263)(530,263)(530,309)(471,309){1}
wire [3:0] w5;    //: /sn:0 {0}(392,157)(392,231)(425,231)(425,280){1}
//: enddecls

  concat g4 (.I0(w3), .I1(w4), .Z(w0));   //: @(357,305) /sn:0 /R:2 /w:[ 1 1 1 ] /dr:0
  //: switch g3 (w1) @(497,263) /sn:0 /w:[ 0 ] /st:0
  //: dip g2 (w6) @(484,146) /sn:0 /w:[ 0 ] /st:7
  //: dip g1 (w5) @(392,147) /sn:0 /w:[ 0 ] /st:7
  led g5 (.I(w0));   //: @(315,229) /sn:0 /w:[ 0 ] /type:3
  CLA g0 (.a(w5), .b(w6), .c_in(w1), .c_out(w4), .s(w3));   //: @(407, 281) /sz:(63, 57) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]

endmodule

module CLA(s, b, c_in, a, c_out);
//: interface  /sz:(63, 57) /bd:[ Ti0>b[3:0](43/63) Ti1>a[3:0](18/63) Ri0>c_in(28/57) Lo0<c_out(29/57) Bo0<s[3:0](31/63) ]
input [3:0] b;    //: /sn:0 {0}(196,40)(236,40){1}
//: {2}(237,40)(307,40){3}
//: {4}(308,40)(379,40){5}
//: {6}(380,40)(450,40){7}
//: {8}(451,40)(558,40){9}
output c_out;    //: /sn:0 {0}(125,222)(200,222){1}
input c_in;    //: /sn:0 /dp:3 {0}(468,107)(500,107){1}
//: {2}(504,107)(557,107){3}
//: {4}(502,109)(502,224)(468,224){5}
output [3:0] s;    //: /sn:0 /dp:1 {0}(166,167)(126,167){1}
input [3:0] a;    //: /sn:0 {0}(196,23)(214,23){1}
//: {2}(215,23)(285,23){3}
//: {4}(286,23)(357,23){5}
//: {6}(358,23)(428,23){7}
//: {8}(429,23)(558,23){9}
wire w13;    //: /sn:0 {0}(451,80)(451,44){1}
wire w6;    //: /sn:0 /dp:1 {0}(226,203)(226,132){1}
wire w7;    //: /sn:0 /dp:1 {0}(210,203)(210,132){1}
wire w25;    //: /sn:0 {0}(308,80)(308,44){1}
wire w4;    //: /sn:0 /dp:1 {0}(297,203)(297,132){1}
wire w36;    //: /sn:0 /dp:1 {0}(172,182)(242,182)(242,132){1}
wire w3;    //: /sn:0 /dp:1 {0}(353,203)(353,132){1}
wire w0;    //: /sn:0 /dp:1 {0}(440,203)(440,132){1}
wire w20;    //: /sn:0 {0}(358,80)(358,27){1}
wire w19;    //: /sn:0 {0}(380,80)(380,44){1}
wire w18;    //: /sn:0 {0}(456,132)(456,152)(172,152){1}
wire w24;    //: /sn:0 {0}(385,132)(385,162)(172,162){1}
wire w31;    //: /sn:0 {0}(237,80)(237,44){1}
wire w1;    //: /sn:0 /dp:1 {0}(424,203)(424,132){1}
wire w32;    //: /sn:0 {0}(215,80)(215,27){1}
wire w27;    //: /sn:0 {0}(325,107)(334,107)(334,203){1}
wire w14;    //: /sn:0 {0}(429,80)(429,27){1}
wire w11;    //: /sn:0 /dp:1 {0}(263,203)(263,107)(254,107){1}
wire w2;    //: /sn:0 /dp:1 {0}(369,203)(369,132){1}
wire w15;    //: /sn:0 {0}(172,172)(313,172)(313,132){1}
wire w5;    //: /sn:0 /dp:1 {0}(281,203)(281,132){1}
wire w26;    //: /sn:0 {0}(286,80)(286,27){1}
wire w9;    //: /sn:0 /dp:1 {0}(405,203)(405,107)(397,107){1}
//: enddecls

  //: joint g8 (c_in) @(502, 107) /w:[ 2 -1 1 4 ]
  PFA g4 (.a(w32), .b(w31), .c(w11), .s(w36), .g(w6), .p(w7));   //: @(201, 81) /sz:(52, 50) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Bo0<1 Bo1<1 Bo2<1 ]
  tran g16(.Z(w32), .I(a[3]));   //: @(215,21) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  PFA g3 (.a(w26), .b(w25), .c(w27), .s(w15), .g(w4), .p(w5));   //: @(272, 81) /sz:(52, 50) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>0 Bo0<1 Bo1<1 Bo2<1 ]
  //: output g17 (s) @(129,167) /sn:0 /R:2 /w:[ 1 ]
  PFA g2 (.a(w20), .b(w19), .c(w9), .s(w24), .g(w2), .p(w3));   //: @(344, 81) /sz:(52, 50) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Bo0<0 Bo1<1 Bo2<1 ]
  PFA g1 (.a(w14), .b(w13), .c(c_in), .s(w18), .g(w0), .p(w1));   //: @(415, 81) /sz:(52, 50) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>0 Bo0<0 Bo1<1 Bo2<1 ]
  concat g18 (.I0(w18), .I1(w24), .I2(w15), .I3(w36), .Z(s));   //: @(167,167) /sn:0 /R:2 /w:[ 1 1 0 0 0 ] /dr:0
  tran g10(.Z(w19), .I(b[1]));   //: @(380,38) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  //: input g6 (b) @(560,40) /sn:0 /R:2 /w:[ 9 ]
  tran g9(.Z(w13), .I(b[0]));   //: @(451,38) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  //: input g7 (c_in) @(559,107) /sn:0 /R:2 /w:[ 3 ]
  tran g12(.Z(w31), .I(b[3]));   //: @(237,38) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  tran g14(.Z(w20), .I(a[1]));   //: @(358,21) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  tran g11(.Z(w25), .I(b[2]));   //: @(308,38) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  //: input g5 (a) @(560,23) /sn:0 /R:2 /w:[ 9 ]
  //: output g19 (c_out) @(128,222) /sn:0 /R:2 /w:[ 0 ]
  tran g15(.Z(w26), .I(a[2]));   //: @(286,21) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  CarryLookaheadLogic g0 (.p3(w7), .g3(w6), .p2(w5), .g2(w4), .p1(w3), .g1(w2), .p0(w1), .g0(w0), .c0(c_in), .c3(w11), .c2(w27), .c1(w9), .c4(c_out));   //: @(201, 204) /sz:(266, 40) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>0 Ti3>0 Ti4>0 Ti5>0 Ti6>0 Ti7>0 Ri0>5 To0<0 To1<1 To2<0 Lo0<1 ]
  tran g13(.Z(w14), .I(a[0]));   //: @(429,21) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1

endmodule
