//: version "1.8.7"

module CSA(c_in, b, a, c_out, s);
//: interface  /sz:(129, 81) /bd:[ Ti0>a[3:0](31/129) Ti1>b[3:0](86/129) Ri0>c_in(40/81) Lo0<c_out(38/81) Bo0<s[3:0](65/129) ]
input [3:0] b;    //: /sn:0 /dp:3 {0}(327,253)(327,230)(456,230)(456,45){1}
//: {2}(458,43)(581,43){3}
//: {4}(454,43)(328,43)(328,90){5}
output c_out;    //: /sn:0 {0}(11,213)(93,213){1}
input c_in;    //: /sn:0 /dp:3 {0}(106,190)(106,67)(480,67){1}
//: {2}(484,67)(580,67){3}
//: {4}(482,69)(482,398)(168,398)(168,379){5}
output [3:0] s;    //: /sn:0 {0}(11,256)(80,256)(80,356)(155,356){1}
input [3:0] a;    //: /sn:0 /dp:3 {0}(284,253)(284,206)(431,206)(431,18){1}
//: {2}(433,16)(581,16){3}
//: {4}(429,16)(285,16)(285,90){5}
wire w13;    //: /sn:0 /dp:1 {0}(122,223)(154,223)(154,295)(259,295){1}
wire w7;    //: /sn:0 {0}(351,294)(418,294)(418,268)(399,268){1}
wire [3:0] w4;    //: /sn:0 {0}(307,171)(307,192)(193,192)(193,346)(184,346){1}
wire w3;    //: /sn:0 {0}(260,132)(155,132)(155,203)(122,203){1}
wire w2;    //: /sn:0 {0}(352,131)(417,131)(417,105)(396,105){1}
wire [3:0] w9;    //: /sn:0 {0}(306,334)(306,366)(184,366){1}
//: enddecls

  //: joint g8 (a) @(431, 16) /w:[ 2 -1 4 1 ]
  //: input g4 (c_in) @(582,67) /sn:0 /R:2 /w:[ 3 ]
  //: input g3 (b) @(583,43) /sn:0 /R:2 /w:[ 3 ]
  //: input g2 (a) @(583,16) /sn:0 /R:2 /w:[ 3 ]
  CPA g1 (.a(a), .b(b), .c_in(w7), .c_out(w13), .s(w9));   //: @(260, 254) /sz:(90, 79) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>0 Lo0<1 Bo0<0 ]
  mux g10 (.I0(w3), .I1(w13), .S(c_in), .Z(c_out));   //: @(106,213) /sn:0 /R:3 /delay:" 6 6" /w:[ 1 0 0 1 ] /ss:0 /do:0
  //: switch g6 (w7) @(382,268) /sn:0 /w:[ 1 ] /st:1
  //: joint g7 (c_in) @(482, 67) /w:[ 2 -1 1 4 ]
  mux g9 (.I0(w4), .I1(w9), .S(c_in), .Z(s));   //: @(168,356) /sn:0 /R:3 /delay:" 6 6" /w:[ 1 1 5 1 ] /ss:1 /do:0
  //: output g12 (c_out) @(14,213) /sn:0 /R:2 /w:[ 0 ]
  //: joint g11 (b) @(456, 43) /w:[ 2 -1 4 1 ]
  //: switch g5 (w2) @(379,105) /sn:0 /w:[ 1 ] /st:0
  //: frame g14 @(-39,-17) /sn:0 /wi:659 /ht:435 /tx:""
  CPA g0 (.a(a), .b(b), .c_in(w2), .c_out(w3), .s(w4));   //: @(261, 91) /sz:(90, 79) /sn:0 /p:[ Ti0>5 Ti1>5 Ri0>0 Lo0<0 Bo0<0 ]
  //: comment g15 /dolink:0 /link:"" @(-36,-43) /sn:0 /R:2
  //: /line:"Carry Select Adder 4bits"
  //: /end
  //: output g13 (s) @(14,256) /sn:0 /R:2 /w:[ 0 ]

endmodule

module CPA(c_out, s, c_in, b, a);
//: interface  /sz:(90, 79) /bd:[ Ti0>b[3:0](67/90) Ti1>a[3:0](24/90) Ri0>c_in(40/79) Lo0<c_out(41/79) Bo0<s[3:0](46/90) ]
input [3:0] b;    //: /sn:0 {0}(507,173)(428,173){1}
//: {2}(427,173)(342,173){3}
//: {4}(341,173)(257,173){5}
//: {6}(256,173)(170,173){7}
//: {8}(169,173)(157,173){9}
output c_out;    //: /sn:0 /dp:1 {0}(148,269)(53,269){1}
input c_in;    //: /sn:0 {0}(507,212)(476,212)(476,269)(465,269){1}
output [3:0] s;    //: /sn:0 /dp:1 {0}(100,323)(85,323)(85,287)(52,287){1}
input [3:0] a;    //: /sn:0 {0}(507,191)(448,191){1}
//: {2}(447,191)(362,191){3}
//: {4}(361,191)(277,191){5}
//: {6}(276,191)(190,191){7}
//: {8}(189,191)(157,191){9}
wire w6;    //: /sn:0 {0}(342,249)(342,177){1}
wire w16;    //: /sn:0 {0}(170,249)(170,177){1}
wire w4;    //: /sn:0 {0}(436,291)(436,308)(106,308){1}
wire w0;    //: /sn:0 {0}(448,249)(448,195){1}
wire w3;    //: /sn:0 {0}(406,269)(379,269){1}
wire w12;    //: /sn:0 {0}(294,269)(320,269){1}
wire w19;    //: /sn:0 {0}(178,291)(178,338)(106,338){1}
wire w10;    //: /sn:0 {0}(277,249)(277,195){1}
wire w1;    //: /sn:0 {0}(428,249)(428,177){1}
wire w17;    //: /sn:0 {0}(207,269)(235,269){1}
wire w14;    //: /sn:0 {0}(265,291)(265,328)(106,328){1}
wire w11;    //: /sn:0 {0}(257,249)(257,177){1}
wire w15;    //: /sn:0 {0}(190,249)(190,195){1}
wire w5;    //: /sn:0 {0}(362,249)(362,195){1}
wire w9;    //: /sn:0 {0}(350,291)(350,318)(106,318){1}
//: enddecls

  //: output g4 (c_out) @(56,269) /sn:0 /R:2 /w:[ 1 ]
  FA g8 (.b(w16), .a(w15), .c_in(w17), .c_out(c_out), .s(w19));   //: @(149, 250) /sz:(57, 40) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>0 Lo0<0 Bo0<0 ]
  //: output g3 (s) @(55,287) /sn:0 /R:2 /w:[ 1 ]
  tran g16(.Z(w11), .I(b[2]));   //: @(257,171) /sn:0 /R:1 /w:[ 1 6 5 ] /ss:1
  tran g17(.Z(w16), .I(b[3]));   //: @(170,171) /sn:0 /R:1 /w:[ 1 8 7 ] /ss:1
  //: input g2 (c_in) @(509,212) /sn:0 /R:2 /w:[ 0 ]
  //: input g1 (b) @(509,173) /sn:0 /R:2 /w:[ 0 ]
  //: frame g18 @(-13,158) /sn:0 /wi:565 /ht:200 /tx:""
  tran g10(.Z(w0), .I(a[0]));   //: @(448,189) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:1
  FA g6 (.b(w6), .a(w5), .c_in(w3), .c_out(w12), .s(w9));   //: @(321, 250) /sz:(57, 40) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<1 Bo0<0 ]
  FA g7 (.b(w11), .a(w10), .c_in(w12), .c_out(w17), .s(w14));   //: @(236, 250) /sz:(57, 40) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>0 Lo0<1 Bo0<0 ]
  concat g9 (.I0(w4), .I1(w9), .I2(w14), .I3(w19), .Z(s));   //: @(101,323) /sn:0 /R:2 /w:[ 1 1 1 1 0 ] /dr:0
  tran g12(.Z(w10), .I(a[2]));   //: @(277,189) /sn:0 /R:1 /w:[ 1 6 5 ] /ss:1
  FA g5 (.b(w1), .a(w0), .c_in(c_in), .c_out(w3), .s(w4));   //: @(407, 250) /sz:(57, 40) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<0 Bo0<0 ]
  tran g11(.Z(w5), .I(a[1]));   //: @(362,189) /sn:0 /R:1 /w:[ 1 4 3 ] /ss:1
  tran g14(.Z(w1), .I(b[0]));   //: @(428,171) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:1
  //: comment g19 /dolink:0 /link:"" @(-10,135) /sn:0 /R:2
  //: /line:"Carry Propagation Adder 4bits"
  //: /end
  //: input g0 (a) @(509,191) /sn:0 /R:2 /w:[ 0 ]
  tran g15(.Z(w6), .I(b[1]));   //: @(342,171) /sn:0 /R:1 /w:[ 1 4 3 ] /ss:1
  tran g13(.Z(w15), .I(a[3]));   //: @(190,189) /sn:0 /R:1 /w:[ 1 8 7 ] /ss:1

endmodule

module FA(c_out, s, c_in, b, a);
//: interface  /sz:(57, 40) /bd:[ Ti0>a(41/57) Ti1>b(21/57) Ri0>c_in(19/40) Lo0<c_out(19/40) Bo0<s(29/57) ]
input b;    //: /sn:0 {0}(193,35)(193,98){1}
//: {2}(195,100)(233,100){3}
//: {4}(193,102)(193,162)(300,162){5}
output c_out;    //: /sn:0 /dp:1 {0}(372,145)(398,145){1}
input c_in;    //: /sn:0 /dp:1 {0}(209,35)(209,116){1}
//: {2}(211,118)(282,118)(282,103)(299,103){3}
//: {4}(209,120)(209,144)(300,144){5}
output s;    //: /sn:0 /dp:1 {0}(320,101)(398,101){1}
input a;    //: /sn:0 {0}(177,35)(177,93){1}
//: {2}(179,95)(233,95){3}
//: {4}(177,97)(177,167)(300,167){5}
wire w14;    //: /sn:0 {0}(321,165)(334,165)(334,147)(351,147){1}
wire w2;    //: /sn:0 {0}(254,98)(265,98){1}
//: {2}(269,98)(299,98){3}
//: {4}(267,100)(267,139)(300,139){5}
wire w11;    //: /sn:0 {0}(321,142)(351,142){1}
//: enddecls

  //: output g4 (c_out) @(395,145) /sn:0 /w:[ 1 ]
  and g8 (.I0(w2), .I1(c_in), .Z(w11));   //: @(311,142) /sn:0 /delay:" 5" /w:[ 5 5 0 ]
  //: output g3 (s) @(395,101) /sn:0 /w:[ 1 ]
  //: input g2 (c_in) @(209,33) /sn:0 /R:3 /w:[ 0 ]
  //: input g1 (b) @(193,33) /sn:0 /R:3 /w:[ 0 ]
  //: joint g10 (a) @(177, 95) /w:[ 2 1 -1 4 ]
  xor g6 (.I0(w2), .I1(c_in), .Z(s));   //: @(310,101) /sn:0 /delay:" 6" /w:[ 3 3 0 ]
  or g7 (.I0(w11), .I1(w14), .Z(c_out));   //: @(362,145) /sn:0 /delay:" 5" /w:[ 1 1 0 ]
  and g9 (.I0(b), .I1(a), .Z(w14));   //: @(311,165) /sn:0 /delay:" 5" /w:[ 5 5 0 ]
  //: joint g12 (b) @(193, 100) /w:[ 2 1 -1 4 ]
  //: joint g11 (w2) @(267, 98) /w:[ 2 -1 1 4 ]
  xor g5 (.I0(a), .I1(b), .Z(w2));   //: @(244,98) /sn:0 /delay:" 6" /w:[ 3 3 0 ]
  //: input g0 (a) @(177,33) /sn:0 /R:3 /w:[ 0 ]
  //: joint g13 (c_in) @(209, 118) /w:[ 2 1 -1 4 ]

endmodule

module main;    //: root_module
wire [4:0] w7;    //: /sn:0 /dp:1 {0}(342,329)(411,329){1}
wire [3:0] w4;    //: /sn:0 {0}(313,264)(313,334)(336,334){1}
wire w3;    //: /sn:0 {0}(247,220)(228,220)(228,324)(336,324){1}
wire [3:0] w0;    //: /sn:0 /dp:1 {0}(271,181)(271,152){1}
wire [3:0] w1;    //: /sn:0 /dp:1 {0}(360,181)(360,150){1}
wire w5;    //: /sn:0 {0}(412,222)(378,222){1}
//: enddecls

  concat g4 (.I0(w4), .I1(w3), .Z(w7));   //: @(341,329) /sn:0 /w:[ 1 1 0 ] /dr:0
  //: switch g3 (w5) @(430,222) /sn:0 /R:2 /w:[ 0 ] /st:0
  //: dip g2 (w1) @(360,140) /sn:0 /w:[ 1 ] /st:15
  //: dip g1 (w0) @(271,142) /sn:0 /w:[ 1 ] /st:0
  led g6 (.I(w7));   //: @(418,329) /sn:0 /R:3 /w:[ 1 ] /type:3
  //: comment g7 /dolink:0 /link:"" @(213,98) /sn:0 /R:2
  //: /line:"Carry Select Adder"
  //: /end
  //: frame g5 @(212,115) /sn:0 /wi:255 /ht:249 /tx:""
  CSA g0 (.b(w1), .a(w0), .c_in(w5), .c_out(w3), .s(w4));   //: @(248, 182) /sz:(129, 81) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<0 Bo0<0 ]

endmodule
