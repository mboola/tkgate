//: version "1.8.7"

module full_adder;    //: root_module
wire w4;    //: /sn:0 {0}(119,129)(119,137)(210,137){1}
wire w3;    //: /sn:0 {0}(179,172)(179,181)(240,181)(240,159){1}
wire w0;    //: /sn:0 {0}(179,42)(252,42)(252,117){1}
wire w1;    //: /sn:0 {0}(318,73)(328,73)(328,137)(269,137){1}
wire w5;    //: /sn:0 {0}(175,90)(232,90)(232,117){1}
//: enddecls

  led g4 (.I(w4));   //: @(119,122) /sn:0 /w:[ 0 ] /type:0
  //: switch g3 (w1) @(301,73) /sn:0 /w:[ 0 ] /st:0
  //: switch g2 (w0) @(162,42) /sn:0 /w:[ 0 ] /st:0
  //: switch g1 (w5) @(158,90) /sn:0 /w:[ 0 ] /st:0
  led g5 (.I(w3));   //: @(179,165) /sn:0 /w:[ 0 ] /type:0
  FA g0 (.a(w0), .b(w5), .c_in(w1), .c_out(w4), .s(w3));   //: @(211, 118) /sz:(57, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<1 Bo0<1 ]

endmodule

module FA(c_out, s, c_in, b, a);
//: interface  /sz:(57, 40) /bd:[ Ti0>b(15/40) Ti1>a(29/40) Ri0>c_in(19/40) Lo0<c_out(19/40) Bo0<s(21/40) ]
input b;    //: /sn:0 {0}(76,79)(115,79){1}
//: {2}(119,79)(135,79){3}
//: {4}(117,81)(117,165)(205,165){5}
output c_out;    //: /sn:0 /dp:1 {0}(308,152)(359,152){1}
input c_in;    //: /sn:0 /dp:1 {0}(269,92)(182,92)(182,109){1}
//: {2}(180,111)(79,111){3}
//: {4}(182,113)(182,135)(203,135){5}
output s;    //: /sn:0 /dp:1 {0}(290,90)(359,90){1}
input a;    //: /sn:0 {0}(75,55)(97,55){1}
//: {2}(101,55)(127,55)(127,74)(135,74){3}
//: {4}(99,57)(99,170)(205,170){5}
wire w14;    //: /sn:0 {0}(226,168)(277,168)(277,154)(287,154){1}
wire w11;    //: /sn:0 {0}(224,138)(277,138)(277,149)(287,149){1}
wire w2;    //: /sn:0 {0}(156,77)(171,77){1}
//: {2}(175,77)(234,77)(234,87)(269,87){3}
//: {4}(173,79)(173,140)(203,140){5}
//: enddecls

  and g8 (.I0(c_in), .I1(w2), .Z(w11));   //: @(214,138) /sn:0 /w:[ 5 5 0 ]
  //: output g4 (c_out) @(356,152) /sn:0 /w:[ 1 ]
  //: output g3 (s) @(356,90) /sn:0 /w:[ 1 ]
  //: input g2 (c_in) @(77,111) /sn:0 /w:[ 3 ]
  //: input g1 (b) @(74,79) /sn:0 /w:[ 0 ]
  //: joint g10 (c_in) @(182, 111) /w:[ -1 1 2 4 ]
  xor g6 (.I0(w2), .I1(c_in), .Z(s));   //: @(280,90) /sn:0 /w:[ 3 0 0 ]
  and g9 (.I0(b), .I1(a), .Z(w14));   //: @(216,168) /sn:0 /w:[ 5 5 0 ]
  or g7 (.I0(w11), .I1(w14), .Z(c_out));   //: @(298,152) /sn:0 /w:[ 1 1 0 ]
  //: joint g12 (b) @(117, 79) /w:[ 2 -1 1 4 ]
  //: joint g11 (w2) @(173, 77) /w:[ 2 -1 1 4 ]
  xor g5 (.I0(a), .I1(b), .Z(w2));   //: @(146,77) /sn:0 /w:[ 3 3 0 ]
  //: input g0 (a) @(73,55) /sn:0 /w:[ 0 ]
  //: joint g13 (a) @(99, 55) /w:[ 2 -1 1 4 ]

endmodule
