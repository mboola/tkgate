//: version "1.8.7"

module CSA(c_in, b, a, c_out, s);
//: interface  /sz:(129, 81) /bd:[ Ti0>a[3:0](31/129) Ti1>b[3:0](86/129) Ri0>c_in(40/81) Lo0<c_out(38/81) Bo0<s[3:0](65/129) ]
input [3:0] b;    //: /sn:0 /dp:3 {0}(733,359)(733,336)(862,336)(862,151){1}
//: {2}(864,149)(987,149){3}
//: {4}(860,149)(734,149)(734,196){5}
output c_out;    //: /sn:0 {0}(417,319)(499,319){1}
input c_in;    //: /sn:0 /dp:3 {0}(512,296)(512,173)(886,173){1}
//: {2}(890,173)(986,173){3}
//: {4}(888,175)(888,504)(574,504)(574,485){5}
output [3:0] s;    //: /sn:0 {0}(417,362)(486,362)(486,462)(561,462){1}
input [3:0] a;    //: /sn:0 /dp:3 {0}(690,359)(690,312)(837,312)(837,124){1}
//: {2}(839,122)(987,122){3}
//: {4}(835,122)(691,122)(691,196){5}
wire w13;    //: /sn:0 /dp:1 {0}(528,329)(560,329)(560,401)(665,401){1}
wire w7;    //: /sn:0 {0}(757,400)(824,400)(824,374)(805,374){1}
wire [3:0] w4;    //: /sn:0 {0}(713,277)(713,298)(599,298)(599,452)(590,452){1}
wire w3;    //: /sn:0 {0}(666,238)(561,238)(561,309)(528,309){1}
wire w2;    //: /sn:0 {0}(758,237)(823,237)(823,211)(802,211){1}
wire [3:0] w9;    //: /sn:0 {0}(712,440)(712,472)(590,472){1}
//: enddecls

  //: joint g8 (a) @(837, 122) /w:[ 2 -1 4 1 ]
  //: input g4 (c_in) @(988,173) /sn:0 /R:2 /w:[ 3 ]
  //: input g3 (b) @(989,149) /sn:0 /R:2 /w:[ 3 ]
  //: input g2 (a) @(989,122) /sn:0 /R:2 /w:[ 3 ]
  CPA g1 (.a(a), .b(b), .c_in(w7), .c_out(w13), .s(w9));   //: @(666, 360) /sz:(90, 79) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>0 Lo0<1 Bo0<0 ]
  mux g10 (.I0(w3), .I1(w13), .S(c_in), .Z(c_out));   //: @(512,319) /sn:0 /R:3 /delay:" 6 6" /w:[ 1 0 0 1 ] /ss:0 /do:0
  //: switch g6 (w7) @(788,374) /sn:0 /w:[ 1 ] /st:1
  //: joint g7 (c_in) @(888, 173) /w:[ 2 -1 1 4 ]
  mux g9 (.I0(w4), .I1(w9), .S(c_in), .Z(s));   //: @(574,462) /sn:0 /R:3 /delay:" 6 6" /w:[ 1 1 5 1 ] /ss:1 /do:0
  //: output g12 (c_out) @(420,319) /sn:0 /R:2 /w:[ 0 ]
  //: joint g11 (b) @(862, 149) /w:[ 2 -1 4 1 ]
  //: switch g5 (w2) @(785,211) /sn:0 /w:[ 1 ] /st:0
  CPA g0 (.a(a), .b(b), .c_in(w2), .c_out(w3), .s(w4));   //: @(667, 197) /sz:(90, 79) /sn:0 /p:[ Ti0>5 Ti1>5 Ri0>0 Lo0<0 Bo0<0 ]
  //: output g13 (s) @(420,362) /sn:0 /R:2 /w:[ 0 ]

endmodule

module CPA(c_out, s, c_in, b, a);
//: interface  /sz:(90, 79) /bd:[ Ti0>b[3:0](67/90) Ti1>a[3:0](24/90) Ri0>c_in(40/79) Lo0<c_out(41/79) Bo0<s[3:0](46/90) ]
input [3:0] b;    //: /sn:0 {0}(507,173)(428,173){1}
//: {2}(427,173)(342,173){3}
//: {4}(341,173)(257,173){5}
//: {6}(256,173)(170,173){7}
//: {8}(169,173)(157,173){9}
output c_out;    //: /sn:0 /dp:1 {0}(148,269)(53,269){1}
input c_in;    //: /sn:0 {0}(507,212)(476,212)(476,269)(465,269){1}
output [3:0] s;    //: /sn:0 /dp:1 {0}(100,323)(85,323)(85,287)(52,287){1}
input [3:0] a;    //: /sn:0 {0}(507,191)(448,191){1}
//: {2}(447,191)(362,191){3}
//: {4}(361,191)(277,191){5}
//: {6}(276,191)(190,191){7}
//: {8}(189,191)(157,191){9}
wire w6;    //: /sn:0 {0}(342,249)(342,177){1}
wire w16;    //: /sn:0 {0}(170,249)(170,177){1}
wire w4;    //: /sn:0 {0}(436,291)(436,308)(106,308){1}
wire w0;    //: /sn:0 {0}(448,249)(448,195){1}
wire w3;    //: /sn:0 {0}(406,269)(379,269){1}
wire w12;    //: /sn:0 {0}(294,269)(320,269){1}
wire w19;    //: /sn:0 {0}(178,291)(178,338)(106,338){1}
wire w10;    //: /sn:0 {0}(277,249)(277,195){1}
wire w1;    //: /sn:0 {0}(428,249)(428,177){1}
wire w17;    //: /sn:0 {0}(207,269)(235,269){1}
wire w14;    //: /sn:0 {0}(265,291)(265,328)(106,328){1}
wire w11;    //: /sn:0 {0}(257,249)(257,177){1}
wire w15;    //: /sn:0 {0}(190,249)(190,195){1}
wire w5;    //: /sn:0 {0}(362,249)(362,195){1}
wire w9;    //: /sn:0 {0}(350,291)(350,318)(106,318){1}
//: enddecls

  //: output g4 (c_out) @(56,269) /sn:0 /R:2 /w:[ 1 ]
  FA g8 (.b(w16), .a(w15), .c_in(w17), .c_out(c_out), .s(w19));   //: @(149, 250) /sz:(57, 40) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>0 Lo0<0 Bo0<0 ]
  //: output g3 (s) @(55,287) /sn:0 /R:2 /w:[ 1 ]
  tran g16(.Z(w11), .I(b[2]));   //: @(257,171) /sn:0 /R:1 /w:[ 1 6 5 ] /ss:1
  tran g17(.Z(w16), .I(b[3]));   //: @(170,171) /sn:0 /R:1 /w:[ 1 8 7 ] /ss:1
  //: input g2 (c_in) @(509,212) /sn:0 /R:2 /w:[ 0 ]
  //: input g1 (b) @(509,173) /sn:0 /R:2 /w:[ 0 ]
  tran g10(.Z(w0), .I(a[0]));   //: @(448,189) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:1
  FA g6 (.b(w6), .a(w5), .c_in(w3), .c_out(w12), .s(w9));   //: @(321, 250) /sz:(57, 40) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<1 Bo0<0 ]
  FA g7 (.b(w11), .a(w10), .c_in(w12), .c_out(w17), .s(w14));   //: @(236, 250) /sz:(57, 40) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>0 Lo0<1 Bo0<0 ]
  concat g9 (.I0(w4), .I1(w9), .I2(w14), .I3(w19), .Z(s));   //: @(101,323) /sn:0 /R:2 /w:[ 1 1 1 1 0 ] /dr:0
  tran g12(.Z(w10), .I(a[2]));   //: @(277,189) /sn:0 /R:1 /w:[ 1 6 5 ] /ss:1
  FA g5 (.b(w1), .a(w0), .c_in(c_in), .c_out(w3), .s(w4));   //: @(407, 250) /sz:(57, 40) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<0 Bo0<0 ]
  tran g11(.Z(w5), .I(a[1]));   //: @(362,189) /sn:0 /R:1 /w:[ 1 4 3 ] /ss:1
  tran g14(.Z(w1), .I(b[0]));   //: @(428,171) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:1
  //: input g0 (a) @(509,191) /sn:0 /R:2 /w:[ 0 ]
  tran g15(.Z(w6), .I(b[1]));   //: @(342,171) /sn:0 /R:1 /w:[ 1 4 3 ] /ss:1
  tran g13(.Z(w15), .I(a[3]));   //: @(190,189) /sn:0 /R:1 /w:[ 1 8 7 ] /ss:1

endmodule

module CSA16(s, c_in, b, c_out, a);
//: interface  /sz:(93, 92) /bd:[ Ti0>b[15:0](29/93) Ti1>a[15:0](63/93) Ri0>c_in(44/92) Lo0<c_out(44/92) Bo0<s[15:0](44/93) ]
input [15:0] b;    //: /sn:0 {0}(603,231)(533,231){1}
//: {2}(532,231)(396,231){3}
//: {4}(395,231)(243,231){5}
//: {6}(242,231)(87,231){7}
//: {8}(86,231)(19,231){9}
output c_out;    //: /sn:0 {0}(-88,357)(0,357){1}
input c_in;    //: /sn:0 /dp:1 {0}(558,360)(580,360)(580,279)(605,279){1}
output [15:0] s;    //: /sn:0 /dp:1 {0}(-27,439)(-52,439)(-52,382)(-87,382){1}
input [15:0] a;    //: /sn:0 {0}(603,255)(489,255){1}
//: {2}(488,255)(341,255){3}
//: {4}(340,255)(188,255){5}
//: {6}(187,255)(32,255){7}
//: {8}(31,255)(18,255){9}
wire [3:0] w6;    //: /sn:0 {0}(396,318)(396,235){1}
wire [3:0] w16;    //: /sn:0 {0}(66,401)(66,424)(-21,424){1}
wire [3:0] w13;    //: /sn:0 {0}(87,318)(87,235){1}
wire [3:0] w7;    //: /sn:0 {0}(32,318)(32,259){1}
wire [3:0] w3;    //: /sn:0 {0}(243,318)(243,235){1}
wire [3:0] w0;    //: /sn:0 {0}(533,318)(533,235){1}
wire [3:0] w12;    //: /sn:0 {0}(222,401)(222,434)(-21,434){1}
wire [3:0] w19;    //: /sn:0 /dp:1 {0}(-21,454)(512,454)(512,401){1}
wire [3:0] w18;    //: /sn:0 /dp:1 {0}(-21,444)(375,444)(375,401){1}
wire [3:0] w1;    //: /sn:0 {0}(489,318)(489,259){1}
wire w8;    //: /sn:0 {0}(440,359)(464,359){1}
wire w14;    //: /sn:0 {0}(131,357)(156,357){1}
wire [3:0] w2;    //: /sn:0 {0}(188,318)(188,259){1}
wire [3:0] w5;    //: /sn:0 {0}(341,318)(341,259){1}
wire w9;    //: /sn:0 {0}(287,358)(309,358){1}
//: enddecls

  CSA g4 (.b(w6), .a(w5), .c_in(w8), .c_out(w9), .s(w18));   //: @(310, 319) /sz:(129, 81) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>0 Lo0<1 Bo0<1 ]
  tran g8(.Z(w1), .I(a[3:0]));   //: @(489,253) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:1
  concat g16 (.I0(w19), .I1(w18), .I2(w12), .I3(w16), .Z(s));   //: @(-26,439) /sn:0 /R:2 /w:[ 0 0 1 1 0 ] /dr:1
  CPA g3 (.a(w1), .b(w0), .c_in(c_in), .c_out(w8), .s(w19));   //: @(465, 319) /sz:(92, 81) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>0 Lo0<1 Bo0<1 ]
  //: output g17 (s) @(-84,382) /sn:0 /R:2 /w:[ 1 ]
  //: input g2 (c_in) @(607,279) /sn:0 /R:2 /w:[ 1 ]
  //: input g1 (b) @(605,231) /sn:0 /R:2 /w:[ 0 ]
  //: frame g18 @(-126,208) /sn:0 /wi:775 /ht:267 /tx:""
  tran g10(.Z(w5), .I(a[7:4]));   //: @(341,253) /sn:0 /R:1 /w:[ 1 4 3 ] /ss:1
  CSA g6 (.b(w13), .a(w7), .c_in(w14), .c_out(c_out), .s(w16));   //: @(1, 319) /sz:(129, 81) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>0 Lo0<1 Bo0<0 ]
  tran g9(.Z(w6), .I(b[7:4]));   //: @(396,229) /sn:0 /R:1 /w:[ 1 4 3 ] /ss:1
  tran g7(.Z(w0), .I(b[3:0]));   //: @(533,229) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:1
  tran g12(.Z(w2), .I(a[11:8]));   //: @(188,253) /sn:0 /R:1 /w:[ 1 6 5 ] /ss:1
  tran g14(.Z(w7), .I(a[15:12]));   //: @(32,253) /sn:0 /R:1 /w:[ 1 8 7 ] /ss:1
  tran g11(.Z(w3), .I(b[11:8]));   //: @(243,229) /sn:0 /R:1 /w:[ 1 6 5 ] /ss:1
  CSA g5 (.b(w3), .a(w2), .c_in(w9), .c_out(w14), .s(w12));   //: @(157, 319) /sz:(129, 81) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>0 Lo0<1 Bo0<0 ]
  //: comment g19 /dolink:0 /link:"" @(-125,184) /sn:0 /R:2
  //: /line:"Carry Select Adder 16bits + Carry Propagate Adder 4bits"
  //: /end
  //: output g15 (c_out) @(-85,357) /sn:0 /R:2 /w:[ 0 ]
  //: input g0 (a) @(605,255) /sn:0 /R:2 /w:[ 0 ]
  tran g13(.Z(w13), .I(b[15:12]));   //: @(87,229) /sn:0 /R:1 /w:[ 1 8 7 ] /ss:1

endmodule

module main;    //: root_module
wire [15:0] w3;    //: /sn:0 /dp:1 {0}(352,168)(352,301)(510,301)(510,289){1}
wire [15:0] w0;    //: /sn:0 /dp:1 {0}(561,115)(561,152)(529,152)(529,195){1}
wire w1;    //: /sn:0 /dp:1 {0}(431,206)(431,240)(465,240){1}
wire [15:0] w2;    //: /sn:0 /dp:1 {0}(495,195)(495,152)(463,152)(463,115){1}
wire w5;    //: /sn:0 {0}(647,105)(627,105)(627,240)(560,240){1}
//: enddecls

  led g4 (.I(w1));   //: @(431,199) /sn:0 /w:[ 0 ] /type:0
  //: dip g3 (w2) @(463,105) /sn:0 /w:[ 1 ] /st:3839
  //: dip g2 (w0) @(561,105) /sn:0 /w:[ 0 ] /st:65535
  //: switch g1 (w5) @(665,105) /sn:0 /R:2 /w:[ 0 ] /st:1
  //: frame g6 @(227,74) /sn:0 /wi:479 /ht:248 /tx:""
  //: comment g7 /dolink:0 /link:"" @(229,51) /sn:0 /R:2
  //: /line:"Carry Select Adder"
  //: /end
  led g5 (.I(w3));   //: @(352,161) /sn:0 /w:[ 0 ] /type:3
  CSA16 g0 (.b(w2), .a(w0), .c_in(w5), .c_out(w1), .s(w3));   //: @(466, 196) /sz:(93, 92) /sn:0 /p:[ Ti0>0 Ti1>1 Ri0>1 Lo0<1 Bo0<1 ]

endmodule

module FA(c_out, s, c_in, b, a);
//: interface  /sz:(57, 40) /bd:[ Ti0>a(41/57) Ti1>b(21/57) Ri0>c_in(19/40) Lo0<c_out(19/40) Bo0<s(29/57) ]
input b;    //: /sn:0 {0}(193,35)(193,98){1}
//: {2}(195,100)(233,100){3}
//: {4}(193,102)(193,162)(300,162){5}
output c_out;    //: /sn:0 /dp:1 {0}(372,145)(398,145){1}
input c_in;    //: /sn:0 /dp:1 {0}(209,35)(209,116){1}
//: {2}(211,118)(282,118)(282,103)(299,103){3}
//: {4}(209,120)(209,144)(300,144){5}
output s;    //: /sn:0 /dp:1 {0}(320,101)(398,101){1}
input a;    //: /sn:0 {0}(177,35)(177,93){1}
//: {2}(179,95)(233,95){3}
//: {4}(177,97)(177,167)(300,167){5}
wire w14;    //: /sn:0 {0}(321,165)(334,165)(334,147)(351,147){1}
wire w2;    //: /sn:0 {0}(254,98)(265,98){1}
//: {2}(269,98)(299,98){3}
//: {4}(267,100)(267,139)(300,139){5}
wire w11;    //: /sn:0 {0}(321,142)(351,142){1}
//: enddecls

  //: output g4 (c_out) @(395,145) /sn:0 /w:[ 1 ]
  and g8 (.I0(w2), .I1(c_in), .Z(w11));   //: @(311,142) /sn:0 /delay:" 5" /w:[ 5 5 0 ]
  //: output g3 (s) @(395,101) /sn:0 /w:[ 1 ]
  //: input g2 (c_in) @(209,33) /sn:0 /R:3 /w:[ 0 ]
  //: input g1 (b) @(193,33) /sn:0 /R:3 /w:[ 0 ]
  //: joint g10 (a) @(177, 95) /w:[ 2 1 -1 4 ]
  xor g6 (.I0(w2), .I1(c_in), .Z(s));   //: @(310,101) /sn:0 /delay:" 6" /w:[ 3 3 0 ]
  or g7 (.I0(w11), .I1(w14), .Z(c_out));   //: @(362,145) /sn:0 /delay:" 5" /w:[ 1 1 0 ]
  and g9 (.I0(b), .I1(a), .Z(w14));   //: @(311,165) /sn:0 /delay:" 5" /w:[ 5 5 0 ]
  //: joint g12 (b) @(193, 100) /w:[ 2 1 -1 4 ]
  //: joint g11 (w2) @(267, 98) /w:[ 2 -1 1 4 ]
  xor g5 (.I0(a), .I1(b), .Z(w2));   //: @(244,98) /sn:0 /delay:" 6" /w:[ 3 3 0 ]
  //: input g0 (a) @(177,33) /sn:0 /R:3 /w:[ 0 ]
  //: joint g13 (c_in) @(209, 118) /w:[ 2 1 -1 4 ]

endmodule
