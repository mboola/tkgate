//: version "1.8.7"

module PFA(p, c, b, g, s, a);
//: interface  /sz:(52, 50) /bd:[ Ti0>a(14/52) Ti1>b(36/52) Ri0>c(26/50) Bo0<s(41/52) Bo1<g(25/52) Bo2<p(9/52) ]
output p;    //: /sn:0 {0}(506,190)(454,190){1}
input b;    //: /sn:0 {0}(265,98)(265,147){1}
//: {2}(267,149)(341,149){3}
//: {4}(265,151)(265,190){5}
//: {6}(267,192)(433,192){7}
//: {8}(265,194)(265,222)(432,222){9}
output s;    //: /sn:0 /dp:1 {0}(453,159)(506,159){1}
input a;    //: /sn:0 {0}(291,98)(291,142){1}
//: {2}(293,144)(341,144){3}
//: {4}(291,146)(291,185){5}
//: {6}(293,187)(433,187){7}
//: {8}(291,189)(291,217)(432,217){9}
output g;    //: /sn:0 {0}(506,220)(453,220){1}
input c;    //: /sn:0 {0}(242,98)(242,161)(432,161){1}
wire w2;    //: /sn:0 {0}(362,147)(393,147)(393,156)(432,156){1}
//: enddecls

  //: output g8 (p) @(503,190) /sn:0 /w:[ 0 ]
  xor g4 (.I0(w2), .I1(c), .Z(s));   //: @(443,159) /sn:0 /delay:" 6" /w:[ 1 1 0 ]
  xor g3 (.I0(a), .I1(b), .Z(w2));   //: @(352,147) /sn:0 /delay:" 6" /w:[ 3 3 0 ]
  //: input g2 (c) @(242,96) /sn:0 /R:3 /w:[ 0 ]
  //: input g1 (b) @(265,96) /sn:0 /R:3 /w:[ 0 ]
  //: joint g10 (a) @(291, 144) /w:[ 2 1 -1 4 ]
  and g6 (.I0(a), .I1(b), .Z(g));   //: @(443,220) /sn:0 /delay:" 5" /w:[ 9 9 1 ]
  //: output g9 (g) @(503,220) /sn:0 /w:[ 0 ]
  //: output g7 (s) @(503,159) /sn:0 /w:[ 1 ]
  //: joint g12 (a) @(291, 187) /w:[ 6 5 -1 8 ]
  //: joint g11 (b) @(265, 192) /w:[ 6 5 -1 8 ]
  or g5 (.I0(a), .I1(b), .Z(p));   //: @(444,190) /sn:0 /delay:" 5" /w:[ 7 7 1 ]
  //: input g0 (a) @(291,96) /sn:0 /R:3 /w:[ 0 ]
  //: joint g13 (b) @(265, 149) /w:[ 2 1 -1 4 ]

endmodule

module CarryLookaheadLogic(g3, p3, gg, g2, g1, g0, c2, c3, p1, p2, c4, pg, p0, c1, c0);
//: interface  /sz:(266, 40) /bd:[ Ti0>p3(9/266) Ti1>g3(25/266) Ti2>p2(80/266) Ti3>g2(96/266) Ti4>p1(152/266) Ti5>g1(168/266) Ti6>p0(223/266) Ti7>g0(239/266) Ri0>c0(20/40) To0<c3(62/266) To1<c2(133/266) To2<c1(204/266) Lo0<c4(18/40) Bo0<gg(241/266) Bo1<pg(223/266) ]
input g3;    //: /sn:0 {0}(183,69)(183,558)(278,558)(278,511)(306,511){1}
input g2;    //: /sn:0 {0}(286,338)(266,338)(266,359)(163,359){1}
//: {2}(161,357)(161,69){3}
//: {4}(161,361)(161,535)(219,535){5}
input g1;    //: /sn:0 {0}(221,348)(142,348){1}
//: {2}(140,346)(140,240){3}
//: {4}(142,238)(253,238)(253,224)(287,224){5}
//: {6}(140,236)(140,69){7}
//: {8}(140,350)(140,506)(219,506){9}
input c0;    //: /sn:0 /dp:11 {0}(221,278)(9,278){1}
//: {2}(7,276)(7,181){3}
//: {4}(9,179)(220,179){5}
//: {6}(7,177)(7,118){7}
//: {8}(9,116)(220,116){9}
//: {10}(7,114)(7,69){11}
//: {12}(7,280)(7,403)(221,403){13}
output c1;    //: /sn:0 {0}(359,128)(308,128){1}
output c4;    //: /sn:0 {0}(362,501)(327,501){1}
output pg;    //: /sn:0 /dp:1 {0}(436,662)(472,662){1}
input p3;    //: /sn:0 {0}(220,464)(90,464){1}
//: {2}(88,462)(88,425){3}
//: {4}(90,423)(221,423){5}
//: {6}(88,421)(88,69){7}
//: {8}(88,466)(88,499){9}
//: {10}(90,501)(219,501){11}
//: {12}(88,503)(88,528){13}
//: {14}(90,530)(219,530){15}
//: {16}(88,532)(88,655)(415,655){17}
input p2;    //: /sn:0 {0}(221,418)(71,418){1}
//: {2}(69,416)(69,345){3}
//: {4}(71,343)(221,343){5}
//: {6}(69,341)(69,321){7}
//: {8}(71,319)(221,319){9}
//: {10}(69,317)(69,295){11}
//: {12}(71,293)(221,293){13}
//: {14}(69,291)(69,69){15}
//: {16}(69,420)(69,457){17}
//: {18}(71,459)(220,459){19}
//: {20}(69,461)(69,494){21}
//: {22}(71,496)(219,496){23}
//: {24}(69,498)(69,660)(415,660){25}
input p1;    //: /sn:0 {0}(415,665)(50,665)(50,456){1}
//: {2}(52,454)(220,454){3}
//: {4}(50,452)(50,415){5}
//: {6}(52,413)(221,413){7}
//: {8}(50,411)(50,316){9}
//: {10}(52,314)(221,314){11}
//: {12}(50,312)(50,290){13}
//: {14}(52,288)(221,288){15}
//: {16}(50,286)(50,218){17}
//: {18}(52,216)(220,216){19}
//: {20}(50,214)(50,191){21}
//: {22}(52,189)(220,189){23}
//: {24}(50,187)(50,69){25}
output c3;    //: /sn:0 {0}(361,330)(307,330){1}
output c2;    //: /sn:0 {0}(359,219)(308,219){1}
input p0;    //: /sn:0 /dp:7 {0}(415,670)(32,670)(32,410){1}
//: {2}(34,408)(221,408){3}
//: {4}(32,406)(32,285){5}
//: {6}(34,283)(221,283){7}
//: {8}(32,281)(32,186){9}
//: {10}(34,184)(220,184){11}
//: {12}(32,182)(32,123){13}
//: {14}(34,121)(220,121){15}
//: {16}(32,119)(32,69){17}
input g0;    //: /sn:0 {0}(221,324)(122,324){1}
//: {2}(120,322)(120,223){3}
//: {4}(122,221)(220,221){5}
//: {6}(120,219)(120,132){7}
//: {8}(122,130)(287,130){9}
//: {10}(120,128)(120,69){11}
//: {12}(120,326)(120,469)(220,469){13}
output gg;    //: /sn:0 {0}(471,624)(434,624){1}
wire w4;    //: /sn:0 /dp:1 {0}(286,328)(256,328)(256,319)(242,319){1}
wire w3;    //: /sn:0 /dp:1 {0}(241,119)(251,119)(251,125)(287,125){1}
wire w0;    //: /sn:0 /dp:1 {0}(287,214)(253,214)(253,184)(241,184){1}
wire w1;    //: /sn:0 /dp:1 {0}(287,219)(241,219){1}
wire w8;    //: /sn:0 /dp:1 {0}(306,496)(259,496)(259,463){1}
//: {2}(261,461)(386,461)(386,622)(413,622){3}
//: {4}(257,461)(241,461){5}
wire w17;    //: /sn:0 {0}(413,632)(249,632)(249,503){1}
//: {2}(251,501)(306,501){3}
//: {4}(247,501)(240,501){5}
wire w2;    //: /sn:0 /dp:1 {0}(286,323)(266,323)(266,285)(242,285){1}
wire w15;    //: /sn:0 {0}(413,627)(261,627)(261,535){1}
//: {2}(261,531)(261,506)(306,506){3}
//: {4}(259,533)(240,533){5}
wire w5;    //: /sn:0 /dp:1 {0}(306,491)(276,491)(276,415){1}
//: {2}(278,413)(398,413)(398,617)(413,617){3}
//: {4}(274,413)(242,413){5}
wire w9;    //: /sn:0 {0}(242,346)(256,346)(256,333)(286,333){1}
//: enddecls

  //: input g4 (g3) @(183,67) /sn:0 /R:3 /w:[ 0 ]
  //: input g8 (p3) @(88,67) /sn:0 /R:3 /w:[ 7 ]
  //: joint g44 (p2) @(69, 418) /w:[ 1 2 -1 16 ]
  //: output g47 (gg) @(468,624) /sn:0 /w:[ 0 ]
  //: input g3 (g2) @(161,67) /sn:0 /R:3 /w:[ 3 ]
  //: joint g16 (c0) @(7, 179) /w:[ 4 6 -1 3 ]
  //: joint g26 (c0) @(7, 278) /w:[ 1 2 -1 12 ]
  //: joint g17 (p0) @(32, 184) /w:[ 10 12 -1 9 ]
  //: input g2 (g1) @(140,67) /sn:0 /R:3 /w:[ 7 ]
  //: joint g23 (g1) @(140, 238) /w:[ 4 6 -1 3 ]
  and g30 (.I0(p1), .I1(p2), .I2(g0), .Z(w4));   //: @(232,319) /sn:0 /delay:" 5" /w:[ 11 9 0 1 ]
  //: input g1 (g0) @(120,67) /sn:0 /R:3 /w:[ 11 ]
  //: output g24 (c2) @(356,219) /sn:0 /w:[ 0 ]
  //: output g39 (c3) @(358,330) /sn:0 /w:[ 0 ]
  //: joint g60 (p3) @(88, 530) /w:[ 14 13 -1 16 ]
  //: joint g29 (p2) @(69, 293) /w:[ 12 14 -1 11 ]
  and g51 (.I0(p2), .I1(p3), .I2(g1), .Z(w17));   //: @(230,501) /sn:0 /delay:" 5" /w:[ 23 11 9 5 ]
  //: joint g18 (p1) @(50, 189) /w:[ 22 24 -1 21 ]
  or g10 (.I0(w3), .I1(g0), .Z(c1));   //: @(298,128) /sn:0 /delay:" 5" /w:[ 1 9 1 ]
  and g25 (.I0(c0), .I1(p0), .I2(p1), .I3(p2), .Z(w2));   //: @(232,285) /sn:0 /delay:" 5" /w:[ 0 7 15 13 1 ]
  //: joint g49 (p3) @(88, 464) /w:[ 1 2 -1 8 ]
  and g50 (.I0(p3), .I1(p2), .I2(p1), .I3(p0), .Z(pg));   //: @(426,662) /sn:0 /w:[ 17 25 0 0 0 ]
  //: input g6 (p1) @(50,67) /sn:0 /R:3 /w:[ 25 ]
  //: joint g56 (w8) @(259, 461) /w:[ 2 -1 4 1 ]
  //: input g7 (p2) @(69,67) /sn:0 /R:3 /w:[ 15 ]
  and g9 (.I0(c0), .I1(p0), .Z(w3));   //: @(231,119) /sn:0 /delay:" 5" /w:[ 9 15 0 ]
  //: joint g35 (p2) @(69, 343) /w:[ 4 6 -1 3 ]
  or g58 (.I0(w5), .I1(w8), .I2(w17), .I3(w15), .I4(g3), .Z(c4));   //: @(317,501) /sn:0 /delay:" 5" /w:[ 0 0 3 3 1 1 ]
  //: joint g59 (w17) @(249, 501) /w:[ 2 -1 4 1 ]
  or g22 (.I0(w0), .I1(w1), .I2(g1), .Z(c2));   //: @(298,219) /sn:0 /delay:" 5" /w:[ 0 0 5 1 ]
  //: joint g31 (p1) @(50, 314) /w:[ 10 12 -1 9 ]
  //: joint g54 (w5) @(276, 413) /w:[ 2 -1 4 1 ]
  //: joint g33 (g0) @(120, 324) /w:[ 1 2 -1 12 ]
  //: joint g36 (g1) @(140, 348) /w:[ 1 2 -1 8 ]
  //: joint g45 (p3) @(88, 423) /w:[ 4 6 -1 3 ]
  //: output g41 (c4) @(359,501) /sn:0 /w:[ 0 ]
  or g52 (.I0(w5), .I1(w8), .I2(w15), .I3(w17), .Z(gg));   //: @(424,624) /sn:0 /w:[ 3 3 0 0 1 ]
  //: output g42 (pg) @(469,662) /sn:0 /w:[ 1 ]
  and g40 (.I0(c0), .I1(p0), .I2(p1), .I3(p2), .I4(p3), .Z(w5));   //: @(232,413) /sn:0 /delay:" 5" /w:[ 13 3 7 0 5 5 ]
  //: joint g12 (p0) @(32, 121) /w:[ 14 16 -1 13 ]
  //: joint g57 (w15) @(261, 533) /w:[ -1 2 4 1 ]
  //: joint g28 (p1) @(50, 288) /w:[ 14 16 -1 13 ]
  and g34 (.I0(p2), .I1(g1), .Z(w9));   //: @(232,346) /sn:0 /delay:" 5" /w:[ 5 0 0 ]
  and g46 (.I0(p1), .I1(p2), .I2(p3), .I3(g0), .Z(w8));   //: @(231,461) /sn:0 /delay:" 5" /w:[ 3 19 0 13 5 ]
  //: input g5 (p0) @(32,67) /sn:0 /R:3 /w:[ 17 ]
  //: output g14 (c1) @(356,128) /sn:0 /w:[ 0 ]
  //: joint g11 (c0) @(7, 116) /w:[ 8 10 -1 7 ]
  //: joint g61 (p2) @(69, 496) /w:[ 22 21 -1 24 ]
  and g19 (.I0(p1), .I1(g0), .Z(w1));   //: @(231,219) /sn:0 /delay:" 5" /w:[ 19 5 1 ]
  //: joint g21 (g0) @(120, 221) /w:[ 4 6 -1 3 ]
  //: joint g20 (p1) @(50, 216) /w:[ 18 20 -1 17 ]
  //: joint g32 (p2) @(69, 319) /w:[ 8 10 -1 7 ]
  //: joint g63 (p0) @(32, 408) /w:[ 2 4 -1 1 ]
  //: input g0 (c0) @(7,67) /sn:0 /R:3 /w:[ 11 ]
  and g15 (.I0(c0), .I1(p0), .I2(p1), .Z(w0));   //: @(231,184) /sn:0 /delay:" 5" /w:[ 5 11 23 1 ]
  //: joint g38 (g2) @(161, 359) /w:[ 1 2 -1 4 ]
  //: joint g43 (p1) @(50, 413) /w:[ 6 8 -1 5 ]
  //: joint g27 (p0) @(32, 283) /w:[ 6 8 -1 5 ]
  //: joint g48 (p2) @(69, 459) /w:[ 18 17 -1 20 ]
  //: joint g62 (p1) @(50, 454) /w:[ 2 4 -1 1 ]
  or g37 (.I0(w2), .I1(w4), .I2(w9), .I3(g2), .Z(c3));   //: @(297,330) /sn:0 /delay:" 5" /w:[ 0 0 1 0 1 ]
  and g55 (.I0(p3), .I1(g2), .Z(w15));   //: @(230,533) /sn:0 /delay:" 5" /w:[ 15 5 5 ]
  //: joint g13 (g0) @(120, 130) /w:[ 8 10 -1 7 ]
  //: joint g53 (p3) @(88, 501) /w:[ 10 9 -1 12 ]

endmodule

module CLA16(b, s, a, c_in, gg, c_out, pg);
//: interface  /sz:(53, 50) /bd:[ Ti0>a[15:0](11/63) Ti1>b[15:0](27/53) Ri0>c(29/58) Lo0<c_out(24/50) Bo0<pg(30/53) Bo1<gg(40/53) Bo2<s[15:0](10/53) ]
input [15:0] b;    //: /sn:0 {0}(435,15)(325,15){1}
//: {2}(324,15)(254,15){3}
//: {4}(253,15)(182,15){5}
//: {6}(181,15)(111,15){7}
//: {8}(110,15)(77,15){9}
output pg;    //: /sn:0 {0}(-39,241)(300,241)(300,230){1}
output c_out;    //: /sn:0 {0}(-39,207)(76,207){1}
input c_in;    //: /sn:0 {0}(344,209)(390,209)(390,91){1}
//: {2}(390,87)(390,46)(434,46){3}
//: {4}(388,89)(344,89){5}
output [15:0] s;    //: /sn:0 {0}(-39,153)(6,153){1}
input [15:0] a;    //: /sn:0 {0}(435,-11)(306,-11){1}
//: {2}(305,-11)(235,-11){3}
//: {4}(234,-11)(163,-11){5}
//: {6}(162,-11)(92,-11){7}
//: {8}(91,-11)(76,-11){9}
output gg;    //: /sn:0 {0}(-39,263)(318,263)(318,230){1}
wire [3:0] w6;    //: /sn:0 /dp:1 {0}(12,148)(260,148)(260,116){1}
wire w16;    //: /sn:0 {0}(210,188)(210,89)(201,89){1}
wire [3:0] w34;    //: /sn:0 {0}(111,64)(111,19){1}
wire w25;    //: /sn:0 /dp:1 {0}(157,116)(157,188){1}
wire w4;    //: /sn:0 /dp:1 {0}(300,116)(300,188){1}
wire [3:0] w22;    //: /sn:0 {0}(182,64)(182,19){1}
wire [3:0] w0;    //: /sn:0 {0}(306,64)(306,-7){1}
wire w37;    //: /sn:0 /dp:1 {0}(86,116)(86,188){1}
wire [3:0] w21;    //: /sn:0 {0}(163,64)(163,-7){1}
wire w31;    //: /sn:0 /dp:1 {0}(229,116)(229,188){1}
wire [3:0] w1;    //: /sn:0 {0}(325,64)(325,19){1}
wire w32;    //: /sn:0 /dp:1 {0}(245,116)(245,188){1}
wire [3:0] w8;    //: /sn:0 {0}(12,158)(188,158)(188,116){1}
wire [3:0] w27;    //: /sn:0 {0}(235,64)(235,-7){1}
wire w17;    //: /sn:0 {0}(281,188)(281,89)(273,89){1}
wire [3:0] w33;    //: /sn:0 {0}(92,64)(92,-7){1}
wire [3:0] w28;    //: /sn:0 {0}(254,64)(254,19){1}
wire [3:0] w2;    //: /sn:0 /dp:1 {0}(12,138)(331,138)(331,116){1}
wire w15;    //: /sn:0 {0}(139,188)(139,89)(130,89){1}
wire w38;    //: /sn:0 /dp:1 {0}(102,116)(102,188){1}
wire w5;    //: /sn:0 /dp:1 {0}(316,116)(316,188){1}
wire [3:0] w9;    //: /sn:0 {0}(12,168)(117,168)(117,116){1}
wire w26;    //: /sn:0 /dp:1 {0}(173,116)(173,188){1}
//: enddecls

  //: input g8 (b) @(437,15) /sn:0 /R:2 /w:[ 0 ]
  CLA g4 (.b(w34), .a(w33), .c_in(w15), .gg(w38), .pg(w37), .s(w9));   //: @(78, 65) /sz:(51, 50) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Bo0<0 Bo1<0 Bo2<1 ]
  tran g16(.Z(w33), .I(a[15:12]));   //: @(92,-13) /sn:0 /R:1 /w:[ 1 8 7 ] /ss:1
  CLA g3 (.b(w28), .a(w27), .c_in(w17), .gg(w32), .pg(w31), .s(w6));   //: @(221, 65) /sz:(51, 50) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Bo0<0 Bo1<0 Bo2<1 ]
  //: output g17 (s) @(-36,153) /sn:0 /R:2 /w:[ 0 ]
  CLA g2 (.b(w22), .a(w21), .c_in(w16), .gg(w26), .pg(w25), .s(w8));   //: @(149, 65) /sz:(51, 50) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Bo0<0 Bo1<0 Bo2<1 ]
  CarryLookaheadLogic g1 (.g0(w5), .p0(w4), .g1(w32), .p1(w31), .g2(w26), .p2(w25), .g3(w38), .p3(w37), .c0(c_in), .c1(w17), .c2(w16), .c3(w15), .c4(c_out), .pg(pg), .gg(gg));   //: @(77, 189) /sz:(266, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Ti3>1 Ti4>1 Ti5>1 Ti6>1 Ti7>1 Ri0>0 To0<0 To1<0 To2<0 Lo0<1 Bo0<1 Bo1<1 ]
  concat g18 (.I0(w2), .I1(w6), .I2(w8), .I3(w9), .Z(s));   //: @(7,153) /sn:0 /R:2 /w:[ 0 0 0 0 1 ] /dr:0
  tran g10(.Z(w0), .I(a[3:0]));   //: @(306,-13) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:1
  //: joint g6 (c_in) @(390, 89) /w:[ -1 2 4 1 ]
  tran g9(.Z(w1), .I(b[3:0]));   //: @(325,13) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:1
  //: input g7 (a) @(437,-11) /sn:0 /R:2 /w:[ 0 ]
  tran g12(.Z(w27), .I(a[7:4]));   //: @(235,-13) /sn:0 /R:1 /w:[ 1 4 3 ] /ss:1
  tran g14(.Z(w21), .I(a[11:8]));   //: @(163,-13) /sn:0 /R:1 /w:[ 1 6 5 ] /ss:1
  tran g11(.Z(w28), .I(b[7:4]));   //: @(254,13) /sn:0 /R:1 /w:[ 1 4 3 ] /ss:1
  //: input g5 (c_in) @(436,46) /sn:0 /R:2 /w:[ 3 ]
  //: output g21 (gg) @(-36,263) /sn:0 /R:2 /w:[ 0 ]
  //: output g19 (c_out) @(-36,207) /sn:0 /R:2 /w:[ 0 ]
  //: output g20 (pg) @(-36,241) /sn:0 /R:2 /w:[ 0 ]
  tran g15(.Z(w34), .I(b[15:12]));   //: @(111,13) /sn:0 /R:1 /w:[ 1 8 7 ] /ss:1
  CLA g0 (.b(w1), .a(w0), .c_in(c_in), .gg(w5), .pg(w4), .s(w2));   //: @(292, 65) /sz:(51, 50) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>5 Bo0<0 Bo1<0 Bo2<1 ]
  tran g13(.Z(w22), .I(b[11:8]));   //: @(182,13) /sn:0 /R:1 /w:[ 1 6 5 ] /ss:1

endmodule

module main;    //: root_module
wire [15:0] w6;    //: /sn:0 {0}(410,345)(410,416)(229,416)(229,350){1}
wire [15:0] w7;    //: /sn:0 {0}(311,170)(311,239)(409,239)(409,293){1}
wire w4;    //: /sn:0 {0}(430,345)(430,419)(492,419)(492,409){1}
wire w3;    //: /sn:0 {0}(399,318)(335,318)(335,285){1}
wire [15:0] w0;    //: /sn:0 {0}(522,180)(522,239)(427,239)(427,293){1}
wire w1;    //: /sn:0 {0}(505,279)(557,279)(557,319)(454,319){1}
wire w5;    //: /sn:0 {0}(440,345)(440,397)(468,397)(468,387){1}
//: enddecls

  led g4 (.I(w3));   //: @(335,278) /sn:0 /w:[ 1 ] /type:0
  //: switch g3 (w1) @(488,279) /sn:0 /w:[ 0 ] /st:0
  //: dip g2 (w0) @(522,170) /sn:0 /w:[ 0 ] /st:7
  //: dip g1 (w7) @(311,160) /sn:0 /w:[ 0 ] /st:7
  led g6 (.I(w5));   //: @(468,380) /sn:0 /w:[ 1 ] /type:0
  led g7 (.I(w4));   //: @(492,402) /sn:0 /w:[ 1 ] /type:0
  led g5 (.I(w6));   //: @(229,343) /sn:0 /w:[ 1 ] /type:3
  CLA16 g0 (.b(w0), .a(w7), .c_in(w1), .c_out(w3), .s(w6), .gg(w5), .pg(w4));   //: @(400, 294) /sz:(53, 50) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 Bo1<0 Bo2<0 ]

endmodule

module CLA(pg, s, b, c_in, a, gg, c_out);
//: interface  /sz:(51, 50) /bd:[ Ti0>a[3:0](18/63) Ti1>b[3:0](35/53) Ri0>c_in(28/57) Bo0<s[3:0](41/53) Bo1<pg(9/53) Bo2<gg(25/53) ]
input [3:0] b;    //: /sn:0 {0}(196,40)(236,40){1}
//: {2}(237,40)(307,40){3}
//: {4}(308,40)(379,40){5}
//: {6}(380,40)(450,40){7}
//: {8}(451,40)(558,40){9}
output pg;    //: /sn:0 {0}(124,259)(424,259)(424,245){1}
output c_out;    //: /sn:0 {0}(125,222)(200,222){1}
input c_in;    //: /sn:0 /dp:1 {0}(468,224)(489,224)(489,109){1}
//: {2}(491,107)(557,107){3}
//: {4}(487,107)(468,107){5}
output [3:0] s;    //: /sn:0 /dp:1 {0}(166,167)(126,167){1}
input [3:0] a;    //: /sn:0 {0}(196,23)(214,23){1}
//: {2}(215,23)(285,23){3}
//: {4}(286,23)(357,23){5}
//: {6}(358,23)(428,23){7}
//: {8}(429,23)(558,23){9}
output gg;    //: /sn:0 {0}(124,274)(442,274)(442,245){1}
wire w16;    //: /sn:0 {0}(297,203)(297,132){1}
wire w13;    //: /sn:0 {0}(451,80)(451,44){1}
wire w25;    //: /sn:0 {0}(308,80)(308,44){1}
wire w22;    //: /sn:0 {0}(424,203)(424,132){1}
wire w36;    //: /sn:0 /dp:1 {0}(172,182)(242,182)(242,132){1}
wire w20;    //: /sn:0 {0}(358,80)(358,27){1}
wire w30;    //: /sn:0 {0}(334,203)(334,107)(325,107){1}
wire w29;    //: /sn:0 {0}(263,203)(263,107)(254,107){1}
wire w12;    //: /sn:0 {0}(281,203)(281,132){1}
wire w18;    //: /sn:0 {0}(456,132)(456,152)(172,152){1}
wire w19;    //: /sn:0 {0}(380,80)(380,44){1}
wire w23;    //: /sn:0 {0}(440,203)(440,132){1}
wire w10;    //: /sn:0 {0}(226,203)(226,132){1}
wire w21;    //: /sn:0 {0}(369,203)(369,132){1}
wire w24;    //: /sn:0 {0}(385,132)(385,162)(172,162){1}
wire w31;    //: /sn:0 {0}(237,80)(237,44){1}
wire w32;    //: /sn:0 {0}(215,80)(215,27){1}
wire w8;    //: /sn:0 {0}(210,203)(210,132){1}
wire w17;    //: /sn:0 {0}(353,203)(353,132){1}
wire w33;    //: /sn:0 {0}(405,203)(405,107)(397,107){1}
wire w14;    //: /sn:0 {0}(429,80)(429,27){1}
wire w15;    //: /sn:0 {0}(172,172)(313,172)(313,132){1}
wire w26;    //: /sn:0 {0}(286,80)(286,27){1}
//: enddecls

  //: output g8 (pg) @(127,259) /sn:0 /R:2 /w:[ 0 ]
  PFA g4 (.a(w32), .b(w31), .c(w29), .s(w36), .g(w10), .p(w8));   //: @(201, 81) /sz:(52, 50) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Bo0<1 Bo1<1 Bo2<1 ]
  PFA g3 (.a(w26), .b(w25), .c(w30), .s(w15), .g(w16), .p(w12));   //: @(272, 81) /sz:(52, 50) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Bo0<1 Bo1<1 Bo2<1 ]
  tran g16(.Z(w32), .I(a[3]));   //: @(215,21) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  //: output g17 (s) @(129,167) /sn:0 /R:2 /w:[ 1 ]
  PFA g2 (.a(w20), .b(w19), .c(w33), .s(w24), .g(w21), .p(w17));   //: @(344, 81) /sz:(52, 50) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Bo0<0 Bo1<1 Bo2<1 ]
  PFA g1 (.a(w14), .b(w13), .c(c_in), .s(w18), .g(w23), .p(w22));   //: @(415, 81) /sz:(52, 50) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>5 Bo0<0 Bo1<1 Bo2<1 ]
  concat g18 (.I0(w18), .I1(w24), .I2(w15), .I3(w36), .Z(s));   //: @(167,167) /sn:0 /R:2 /w:[ 1 1 0 0 0 ] /dr:0
  tran g10(.Z(w19), .I(b[1]));   //: @(380,38) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  //: input g6 (b) @(560,40) /sn:0 /R:2 /w:[ 9 ]
  //: input g7 (c_in) @(559,107) /sn:0 /R:2 /w:[ 3 ]
  tran g9(.Z(w13), .I(b[0]));   //: @(451,38) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  tran g12(.Z(w31), .I(b[3]));   //: @(237,38) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  //: input g5 (a) @(560,23) /sn:0 /R:2 /w:[ 9 ]
  tran g11(.Z(w25), .I(b[2]));   //: @(308,38) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  tran g14(.Z(w20), .I(a[1]));   //: @(358,21) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  //: output g21 (gg) @(127,274) /sn:0 /R:2 /w:[ 0 ]
  //: output g19 (c_out) @(128,222) /sn:0 /R:2 /w:[ 0 ]
  CarryLookaheadLogic g20 (.g0(w23), .p0(w22), .g1(w21), .p1(w17), .g2(w16), .p2(w12), .g3(w10), .p3(w8), .c0(c_in), .c1(w33), .c2(w30), .c3(w29), .c4(c_out), .pg(pg), .gg(gg));   //: @(201, 204) /sz:(266, 40) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>0 Ti3>0 Ti4>0 Ti5>0 Ti6>0 Ti7>0 Ri0>0 To0<0 To1<0 To2<0 Lo0<1 Bo0<1 Bo1<1 ]
  //: joint g0 (c_in) @(489, 107) /w:[ 2 -1 4 1 ]
  tran g15(.Z(w26), .I(a[2]));   //: @(286,21) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  tran g13(.Z(w14), .I(a[0]));   //: @(429,21) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1

endmodule
