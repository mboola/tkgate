//: version "1.8.7"

module PFA(p, c, b, g, s, a);
//: interface  /sz:(52, 50) /bd:[ Ti0>a(14/52) Ti1>b(36/52) Ri0>c(26/50) Bo0<s(41/52) Bo1<g(25/52) Bo2<p(9/52) ]
output p;    //: /sn:0 {0}(809,364)(757,364){1}
input b;    //: /sn:0 {0}(568,272)(568,321){1}
//: {2}(570,323)(644,323){3}
//: {4}(568,325)(568,364){5}
//: {6}(570,366)(736,366){7}
//: {8}(568,368)(568,396)(735,396){9}
output s;    //: /sn:0 /dp:1 {0}(756,333)(809,333){1}
input a;    //: /sn:0 {0}(594,272)(594,316){1}
//: {2}(596,318)(644,318){3}
//: {4}(594,320)(594,359){5}
//: {6}(596,361)(736,361){7}
//: {8}(594,363)(594,391)(735,391){9}
output g;    //: /sn:0 {0}(809,394)(756,394){1}
input c;    //: /sn:0 {0}(545,272)(545,335)(735,335){1}
wire w2;    //: /sn:0 {0}(665,321)(696,321)(696,330)(735,330){1}
//: enddecls

  //: output g8 (p) @(806,364) /sn:0 /w:[ 0 ]
  xor g4 (.I0(w2), .I1(c), .Z(s));   //: @(746,333) /sn:0 /delay:" 6" /w:[ 1 1 0 ]
  xor g3 (.I0(a), .I1(b), .Z(w2));   //: @(655,321) /sn:0 /delay:" 6" /w:[ 3 3 0 ]
  //: comment g16 /dolink:0 /link:"" @(826,357) /sn:0
  //: /line:"(T_pn = 5T)"
  //: /end
  //: comment g17 /dolink:0 /link:"" @(825,324) /sn:0
  //: /line:"(T_sn = 12T)"
  //: /end
  //: input g2 (c) @(545,270) /sn:0 /R:3 /w:[ 0 ]
  //: input g1 (b) @(568,270) /sn:0 /R:3 /w:[ 0 ]
  //: comment g18 /dolink:0 /link:"" @(827,384) /sn:0
  //: /line:"(T_gn = 5T)"
  //: /end
  //: joint g10 (a) @(594, 318) /w:[ 2 1 -1 4 ]
  and g6 (.I0(a), .I1(b), .Z(g));   //: @(746,394) /sn:0 /delay:" 5" /w:[ 9 9 1 ]
  //: output g9 (g) @(806,394) /sn:0 /w:[ 0 ]
  //: output g7 (s) @(806,333) /sn:0 /w:[ 1 ]
  //: comment g22 /dolink:0 /link:"" @(742,385) /sn:0
  //: /line:"5T"
  //: /end
  //: joint g12 (a) @(594, 361) /w:[ 6 5 -1 8 ]
  //: joint g11 (b) @(568, 366) /w:[ 6 5 -1 8 ]
  or g5 (.I0(a), .I1(b), .Z(p));   //: @(747,364) /sn:0 /delay:" 5" /w:[ 7 7 1 ]
  //: frame g14 @(522,236) /sn:0 /wi:352 /ht:174 /tx:""
  //: comment g19 /dolink:0 /link:"" @(654,312) /sn:0
  //: /line:"6T"
  //: /end
  //: comment g21 /dolink:0 /link:"" @(744,356) /sn:0
  //: /line:"5T"
  //: /end
  //: comment g20 /dolink:0 /link:"" @(745,324) /sn:0
  //: /line:"6T"
  //: /end
  //: input g0 (a) @(594,270) /sn:0 /R:3 /w:[ 0 ]
  //: comment g15 /dolink:0 /link:"" @(523,217) /sn:0
  //: /line:"Partial Full Adder - Circuit"
  //: /end
  //: joint g13 (b) @(568, 323) /w:[ 2 1 -1 4 ]

endmodule

module CarryLookaheadLogic(g3, p3, gg, g2, g1, g0, c2, c3, p1, p2, c4, pg, p0, c1, c0);
//: interface  /sz:(266, 40) /bd:[ Ti0>p3(9/266) Ti1>g3(25/266) Ti2>p2(80/266) Ti3>g2(96/266) Ti4>p1(152/266) Ti5>g1(168/266) Ti6>p0(223/266) Ti7>g0(239/266) Ri0>c0(20/40) To0<c3(62/266) To1<c2(133/266) To2<c1(204/266) Lo0<c4(18/40) Bo0<gg(241/266) Bo1<pg(223/266) ]
input g3;    //: /sn:0 {0}(183,69)(183,556){1}
//: {2}(185,558)(280,558)(280,511)(306,511){3}
//: {4}(183,560)(183,636)(307,636){5}
input g2;    //: /sn:0 {0}(286,338)(266,338)(266,359)(163,359){1}
//: {2}(161,357)(161,69){3}
//: {4}(161,361)(161,533){5}
//: {6}(163,535)(219,535){7}
//: {8}(161,537)(161,677)(227,677){9}
input g1;    //: /sn:0 {0}(221,348)(142,348){1}
//: {2}(140,346)(140,240){3}
//: {4}(142,238)(254,238)(254,224)(288,224){5}
//: {6}(140,236)(140,69){7}
//: {8}(140,350)(140,506)(219,506){9}
input c0;    //: /sn:0 /dp:11 {0}(221,278)(9,278){1}
//: {2}(7,276)(7,181){3}
//: {4}(9,179)(220,179){5}
//: {6}(7,177)(7,118){7}
//: {8}(9,116)(220,116){9}
//: {10}(7,114)(7,69){11}
//: {12}(7,280)(7,403)(221,403){13}
output c1;    //: /sn:0 {0}(359,128)(308,128){1}
output c4;    //: /sn:0 {0}(362,501)(327,501){1}
input p3;    //: /sn:0 {0}(220,464)(90,464){1}
//: {2}(88,462)(88,425){3}
//: {4}(90,423)(221,423){5}
//: {6}(88,421)(88,69){7}
//: {8}(88,466)(88,499){9}
//: {10}(90,501)(219,501){11}
//: {12}(88,503)(88,528){13}
//: {14}(90,530)(219,530){15}
//: {16}(88,532)(88,575){17}
//: {18}(90,577)(308,577){19}
//: {20}(88,579)(88,603){21}
//: {22}(90,605)(225,605){23}
//: {24}(88,607)(88,641)(225,641){25}
output pg;    //: /sn:0 {0}(377,584)(329,584){1}
input p2;    //: /sn:0 {0}(308,582)(71,582){1}
//: {2}(69,580)(69,498){3}
//: {4}(71,496)(219,496){5}
//: {6}(69,494)(69,461){7}
//: {8}(71,459)(220,459){9}
//: {10}(69,457)(69,420){11}
//: {12}(71,418)(221,418){13}
//: {14}(69,416)(69,345){15}
//: {16}(71,343)(221,343){17}
//: {18}(69,341)(69,321){19}
//: {20}(71,319)(221,319){21}
//: {22}(69,317)(69,295){23}
//: {24}(71,293)(221,293){25}
//: {26}(69,291)(69,69){27}
//: {28}(69,584)(69,608){29}
//: {30}(71,610)(225,610){31}
//: {32}(69,612)(69,644){33}
//: {34}(71,646)(225,646){35}
//: {36}(69,648)(69,672)(227,672){37}
input p1;    //: /sn:0 {0}(225,615)(50,615)(50,589){1}
//: {2}(52,587)(308,587){3}
//: {4}(50,585)(50,456){5}
//: {6}(52,454)(220,454){7}
//: {8}(50,452)(50,415){9}
//: {10}(52,413)(221,413){11}
//: {12}(50,411)(50,316){13}
//: {14}(52,314)(221,314){15}
//: {16}(50,312)(50,290){17}
//: {18}(52,288)(221,288){19}
//: {20}(50,286)(50,218){21}
//: {22}(52,216)(220,216){23}
//: {24}(50,214)(50,191){25}
//: {26}(52,189)(220,189){27}
//: {28}(50,187)(50,69){29}
output c3;    //: /sn:0 {0}(361,330)(307,330){1}
output c2;    //: /sn:0 {0}(359,219)(309,219){1}
input p0;    //: /sn:0 /dp:15 {0}(221,408)(34,408){1}
//: {2}(32,406)(32,285){3}
//: {4}(34,283)(221,283){5}
//: {6}(32,281)(32,186){7}
//: {8}(34,184)(220,184){9}
//: {10}(32,182)(32,123){11}
//: {12}(34,121)(220,121){13}
//: {14}(32,119)(32,69){15}
//: {16}(32,410)(32,592)(308,592){17}
input g0;    //: /sn:0 {0}(225,651)(120,651)(120,622){1}
//: {2}(122,620)(225,620){3}
//: {4}(120,618)(120,471){5}
//: {6}(122,469)(220,469){7}
//: {8}(120,467)(120,326){9}
//: {10}(122,324)(221,324){11}
//: {12}(120,322)(120,223){13}
//: {14}(122,221)(220,221){15}
//: {16}(120,219)(120,132){17}
//: {18}(122,130)(287,130){19}
//: {20}(120,128)(120,69){21}
output gg;    //: /sn:0 /dp:1 {0}(328,643)(374,643){1}
wire w6;    //: /sn:0 {0}(240,501)(306,501){1}
wire w13;    //: /sn:0 /dp:1 {0}(307,651)(293,651)(293,675)(248,675){1}
wire w4;    //: /sn:0 /dp:1 {0}(286,328)(256,328)(256,319)(242,319){1}
wire w3;    //: /sn:0 /dp:1 {0}(241,119)(251,119)(251,125)(287,125){1}
wire w0;    //: /sn:0 /dp:1 {0}(288,214)(254,214)(254,184)(241,184){1}
wire w18;    //: /sn:0 {0}(246,646)(307,646){1}
wire w1;    //: /sn:0 /dp:1 {0}(288,219)(241,219){1}
wire w8;    //: /sn:0 /dp:1 {0}(306,496)(259,496)(259,461)(241,461){1}
wire w14;    //: /sn:0 {0}(246,612)(293,612)(293,641)(307,641){1}
wire w2;    //: /sn:0 /dp:1 {0}(286,323)(266,323)(266,285)(242,285){1}
wire w11;    //: /sn:0 {0}(240,533)(261,533)(261,506)(306,506){1}
wire w5;    //: /sn:0 /dp:1 {0}(306,491)(276,491)(276,413)(242,413){1}
wire w9;    //: /sn:0 {0}(242,346)(256,346)(256,333)(286,333){1}
//: enddecls

  //: input g4 (g3) @(183,67) /sn:0 /R:3 /w:[ 0 ]
  //: input g8 (p3) @(88,67) /sn:0 /R:3 /w:[ 7 ]
  //: joint g44 (p2) @(69, 418) /w:[ 12 14 -1 11 ]
  //: output g47 (gg) @(371,643) /sn:0 /w:[ 1 ]
  //: input g3 (g2) @(161,67) /sn:0 /R:3 /w:[ 3 ]
  //: joint g16 (c0) @(7, 179) /w:[ 4 6 -1 3 ]
  //: joint g26 (c0) @(7, 278) /w:[ 1 2 -1 12 ]
  //: joint g17 (p0) @(32, 184) /w:[ 8 10 -1 7 ]
  //: input g2 (g1) @(140,67) /sn:0 /R:3 /w:[ 7 ]
  //: joint g23 (g1) @(140, 238) /w:[ 4 6 -1 3 ]
  and g30 (.I0(p1), .I1(p2), .I2(g0), .Z(w4));   //: @(232,319) /sn:0 /delay:" 5" /w:[ 15 21 11 1 ]
  //: joint g74 (g3) @(183, 558) /w:[ 2 1 -1 4 ]
  //: input g1 (g0) @(120,67) /sn:0 /R:3 /w:[ 21 ]
  //: output g24 (c2) @(356,219) /sn:0 /w:[ 0 ]
  //: output g39 (c3) @(358,330) /sn:0 /w:[ 0 ]
  //: joint g60 (p3) @(88, 530) /w:[ 14 13 -1 16 ]
  //: joint g29 (p2) @(69, 293) /w:[ 24 26 -1 23 ]
  and g51 (.I0(p2), .I1(p3), .I2(g1), .Z(w6));   //: @(230,501) /sn:0 /delay:" 5" /w:[ 5 11 9 0 ]
  //: joint g18 (p1) @(50, 189) /w:[ 26 28 -1 25 ]
  //: joint g70 (p2) @(69, 610) /w:[ 30 29 -1 32 ]
  or g10 (.I0(w3), .I1(g0), .Z(c1));   //: @(298,128) /sn:0 /delay:" 5" /w:[ 1 19 1 ]
  and g25 (.I0(c0), .I1(p0), .I2(p1), .I3(p2), .Z(w2));   //: @(232,285) /sn:0 /delay:" 5" /w:[ 0 5 19 25 1 ]
  //: frame g65 @(-13,50) /sn:0 /wi:513 /ht:640 /tx:""
  //: comment g64 /dolink:0 /link:"" @(-13,17) /sn:0 /R:2
  //: /line:"Carry Look-Ahead Adder Logic - Circuit"
  //: /end
  //: joint g49 (p3) @(88, 464) /w:[ 1 2 -1 8 ]
  //: joint g72 (p2) @(69, 646) /w:[ 34 33 -1 36 ]
  and g50 (.I0(p3), .I1(p2), .I2(p1), .I3(p0), .Z(pg));   //: @(319,584) /sn:0 /delay:" 5" /w:[ 19 0 3 17 1 ]
  //: input g6 (p1) @(50,67) /sn:0 /R:3 /w:[ 29 ]
  //: input g7 (p2) @(69,67) /sn:0 /R:3 /w:[ 27 ]
  and g9 (.I0(c0), .I1(p0), .Z(w3));   //: @(231,119) /sn:0 /delay:" 5" /w:[ 9 13 0 ]
  //: joint g35 (p2) @(69, 343) /w:[ 16 18 -1 15 ]
  or g58 (.I0(w5), .I1(w8), .I2(w6), .I3(w11), .I4(g3), .Z(c4));   //: @(317,501) /sn:0 /delay:" 5" /w:[ 0 0 1 1 3 1 ]
  //: joint g56 (p3) @(88, 577) /w:[ 18 17 -1 20 ]
  //: joint g68 (g0) @(120, 620) /w:[ 2 4 -1 1 ]
  //: joint g73 (g2) @(161, 535) /w:[ 6 5 -1 8 ]
  or g22 (.I0(w0), .I1(w1), .I2(g1), .Z(c2));   //: @(299,219) /sn:0 /delay:" 5" /w:[ 0 0 5 1 ]
  //: joint g31 (p1) @(50, 314) /w:[ 14 16 -1 13 ]
  //: joint g59 (p1) @(50, 587) /w:[ 2 4 -1 1 ]
  and g71 (.I0(p2), .I1(g2), .Z(w13));   //: @(238,675) /sn:0 /delay:" 5" /w:[ 37 9 1 ]
  and g67 (.I0(p3), .I1(p2), .I2(g0), .Z(w18));   //: @(236,646) /sn:0 /delay:" 5" /w:[ 25 35 0 0 ]
  //: joint g33 (g0) @(120, 324) /w:[ 10 12 -1 9 ]
  //: joint g36 (g1) @(140, 348) /w:[ 1 2 -1 8 ]
  //: joint g45 (p3) @(88, 423) /w:[ 4 6 -1 3 ]
  //: output g41 (c4) @(359,501) /sn:0 /w:[ 0 ]
  and g54 (.I0(p3), .I1(p2), .I2(p1), .I3(g0), .Z(w14));   //: @(236,612) /sn:0 /delay:" 5" /w:[ 23 31 0 3 0 ]
  or g52 (.I0(g3), .I1(w14), .I2(w18), .I3(w13), .Z(gg));   //: @(318,643) /sn:0 /delay:" 5" /w:[ 5 1 1 0 0 ]
  //: output g42 (pg) @(374,584) /sn:0 /w:[ 0 ]
  and g40 (.I0(c0), .I1(p0), .I2(p1), .I3(p2), .I4(p3), .Z(w5));   //: @(232,413) /sn:0 /delay:" 5" /w:[ 13 0 11 13 5 1 ]
  //: joint g69 (p3) @(88, 605) /w:[ 22 21 -1 24 ]
  //: joint g66 (g0) @(120, 469) /w:[ 6 8 -1 5 ]
  //: joint g12 (p0) @(32, 121) /w:[ 12 14 -1 11 ]
  //: joint g28 (p1) @(50, 288) /w:[ 18 20 -1 17 ]
  and g34 (.I0(p2), .I1(g1), .Z(w9));   //: @(232,346) /sn:0 /delay:" 5" /w:[ 17 0 0 ]
  and g46 (.I0(p1), .I1(p2), .I2(p3), .I3(g0), .Z(w8));   //: @(231,461) /sn:0 /delay:" 5" /w:[ 7 9 0 7 1 ]
  //: joint g57 (p2) @(69, 582) /w:[ 1 2 -1 28 ]
  //: input g5 (p0) @(32,67) /sn:0 /R:3 /w:[ 15 ]
  //: output g14 (c1) @(356,128) /sn:0 /w:[ 0 ]
  //: joint g11 (c0) @(7, 116) /w:[ 8 10 -1 7 ]
  //: joint g61 (p2) @(69, 496) /w:[ 4 6 -1 3 ]
  and g19 (.I0(p1), .I1(g0), .Z(w1));   //: @(231,219) /sn:0 /delay:" 5" /w:[ 23 15 1 ]
  //: joint g21 (g0) @(120, 221) /w:[ 14 16 -1 13 ]
  //: joint g20 (p1) @(50, 216) /w:[ 22 24 -1 21 ]
  //: joint g32 (p2) @(69, 319) /w:[ 20 22 -1 19 ]
  //: joint g63 (p0) @(32, 408) /w:[ 1 2 -1 16 ]
  //: input g0 (c0) @(7,67) /sn:0 /R:3 /w:[ 11 ]
  and g15 (.I0(c0), .I1(p0), .I2(p1), .Z(w0));   //: @(231,184) /sn:0 /delay:" 5" /w:[ 5 9 27 1 ]
  //: joint g38 (g2) @(161, 359) /w:[ 1 2 -1 4 ]
  //: joint g43 (p1) @(50, 413) /w:[ 10 12 -1 9 ]
  //: joint g27 (p0) @(32, 283) /w:[ 4 6 -1 3 ]
  //: joint g48 (p2) @(69, 459) /w:[ 8 10 -1 7 ]
  //: joint g62 (p1) @(50, 454) /w:[ 6 8 -1 5 ]
  or g37 (.I0(w2), .I1(w4), .I2(w9), .I3(g2), .Z(c3));   //: @(297,330) /sn:0 /delay:" 5" /w:[ 0 0 1 0 1 ]
  and g55 (.I0(p3), .I1(g2), .Z(w11));   //: @(230,533) /sn:0 /delay:" 5" /w:[ 15 7 0 ]
  //: joint g13 (g0) @(120, 130) /w:[ 18 20 -1 17 ]
  //: joint g53 (p3) @(88, 501) /w:[ 10 9 -1 12 ]

endmodule

module CLA16(b, s, a, c_in, gg, c_out, pg);
//: interface  /sz:(53, 50) /bd:[ Ti0>a[15:0](9/53) Ti1>b[15:0](27/53) Ri0>c(25/50) Lo0<c_out(24/50) Bo0<pg(30/53) Bo1<gg(40/53) Bo2<s[15:0](10/53) ]
input [15:0] b;    //: /sn:0 {0}(435,15)(325,15){1}
//: {2}(324,15)(254,15){3}
//: {4}(253,15)(182,15){5}
//: {6}(181,15)(111,15){7}
//: {8}(110,15)(77,15){9}
output pg;    //: /sn:0 {0}(-39,241)(300,241)(300,230){1}
output c_out;    //: /sn:0 {0}(-39,207)(76,207){1}
input c_in;    //: /sn:0 {0}(344,209)(390,209)(390,91){1}
//: {2}(390,87)(390,46)(434,46){3}
//: {4}(388,89)(344,89){5}
output [15:0] s;    //: /sn:0 {0}(-39,153)(6,153){1}
input [15:0] a;    //: /sn:0 {0}(435,-11)(306,-11){1}
//: {2}(305,-11)(235,-11){3}
//: {4}(234,-11)(163,-11){5}
//: {6}(162,-11)(92,-11){7}
//: {8}(91,-11)(76,-11){9}
output gg;    //: /sn:0 {0}(-39,263)(318,263)(318,230){1}
wire [3:0] w6;    //: /sn:0 /dp:1 {0}(12,148)(260,148)(260,116){1}
wire w16;    //: /sn:0 {0}(210,188)(210,89)(201,89){1}
wire [3:0] w34;    //: /sn:0 {0}(111,64)(111,19){1}
wire w25;    //: /sn:0 /dp:1 {0}(157,116)(157,188){1}
wire w4;    //: /sn:0 /dp:1 {0}(300,116)(300,188){1}
wire [3:0] w22;    //: /sn:0 {0}(182,64)(182,19){1}
wire [3:0] w0;    //: /sn:0 {0}(306,64)(306,-7){1}
wire w37;    //: /sn:0 /dp:1 {0}(86,116)(86,188){1}
wire [3:0] w21;    //: /sn:0 {0}(163,64)(163,-7){1}
wire w31;    //: /sn:0 /dp:1 {0}(229,116)(229,188){1}
wire [3:0] w1;    //: /sn:0 {0}(325,64)(325,19){1}
wire w32;    //: /sn:0 /dp:1 {0}(245,116)(245,188){1}
wire [3:0] w8;    //: /sn:0 {0}(12,158)(188,158)(188,116){1}
wire [3:0] w27;    //: /sn:0 {0}(235,64)(235,-7){1}
wire w17;    //: /sn:0 {0}(281,188)(281,89)(273,89){1}
wire [3:0] w33;    //: /sn:0 {0}(92,64)(92,-7){1}
wire [3:0] w28;    //: /sn:0 {0}(254,64)(254,19){1}
wire [3:0] w2;    //: /sn:0 /dp:1 {0}(12,138)(331,138)(331,116){1}
wire w15;    //: /sn:0 {0}(139,188)(139,89)(130,89){1}
wire w38;    //: /sn:0 /dp:1 {0}(102,116)(102,188){1}
wire w5;    //: /sn:0 /dp:1 {0}(316,116)(316,188){1}
wire [3:0] w9;    //: /sn:0 {0}(12,168)(117,168)(117,116){1}
wire w26;    //: /sn:0 /dp:1 {0}(173,116)(173,188){1}
//: enddecls

  //: input g8 (b) @(437,15) /sn:0 /R:2 /w:[ 0 ]
  CLA g4 (.b(w34), .a(w33), .c_in(w15), .gg(w38), .pg(w37), .s(w9));   //: @(78, 65) /sz:(51, 50) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Bo0<0 Bo1<0 Bo2<1 ]
  tran g16(.Z(w33), .I(a[15:12]));   //: @(92,-13) /sn:0 /R:1 /w:[ 1 8 7 ] /ss:1
  CLA g3 (.b(w28), .a(w27), .c_in(w17), .gg(w32), .pg(w31), .s(w6));   //: @(221, 65) /sz:(51, 50) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Bo0<0 Bo1<0 Bo2<1 ]
  //: output g17 (s) @(-36,153) /sn:0 /R:2 /w:[ 0 ]
  CLA g2 (.b(w22), .a(w21), .c_in(w16), .gg(w26), .pg(w25), .s(w8));   //: @(149, 65) /sz:(51, 50) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Bo0<0 Bo1<0 Bo2<1 ]
  //: comment g23 /dolink:0 /link:"" @(-81,-37) /sn:0 /R:2
  //: /line:"Carry Look-Ahead Adder - Circuit"
  //: /line:""
  //: /end
  CarryLookaheadLogic g1 (.g0(w5), .p0(w4), .g1(w32), .p1(w31), .g2(w26), .p2(w25), .g3(w38), .p3(w37), .c0(c_in), .c1(w17), .c2(w16), .c3(w15), .c4(c_out), .pg(pg), .gg(gg));   //: @(77, 189) /sz:(266, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Ti3>1 Ti4>1 Ti5>1 Ti6>1 Ti7>1 Ri0>0 To0<0 To1<0 To2<0 Lo0<1 Bo0<1 Bo1<1 ]
  concat g18 (.I0(w2), .I1(w6), .I2(w8), .I3(w9), .Z(s));   //: @(7,153) /sn:0 /R:2 /w:[ 0 0 0 0 1 ] /dr:0
  tran g10(.Z(w0), .I(a[3:0]));   //: @(306,-13) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:1
  //: joint g6 (c_in) @(390, 89) /w:[ -1 2 4 1 ]
  tran g9(.Z(w1), .I(b[3:0]));   //: @(325,13) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:1
  //: input g7 (a) @(437,-11) /sn:0 /R:2 /w:[ 0 ]
  //: frame g22 @(-82,-22) /sn:0 /wi:542 /ht:301 /tx:""
  tran g12(.Z(w27), .I(a[7:4]));   //: @(235,-13) /sn:0 /R:1 /w:[ 1 4 3 ] /ss:1
  tran g14(.Z(w21), .I(a[11:8]));   //: @(163,-13) /sn:0 /R:1 /w:[ 1 6 5 ] /ss:1
  tran g11(.Z(w28), .I(b[7:4]));   //: @(254,13) /sn:0 /R:1 /w:[ 1 4 3 ] /ss:1
  //: input g5 (c_in) @(436,46) /sn:0 /R:2 /w:[ 3 ]
  //: output g21 (gg) @(-36,263) /sn:0 /R:2 /w:[ 0 ]
  //: output g19 (c_out) @(-36,207) /sn:0 /R:2 /w:[ 0 ]
  //: output g20 (pg) @(-36,241) /sn:0 /R:2 /w:[ 0 ]
  tran g15(.Z(w34), .I(b[15:12]));   //: @(111,13) /sn:0 /R:1 /w:[ 1 8 7 ] /ss:1
  CLA g0 (.b(w1), .a(w0), .c_in(c_in), .gg(w5), .pg(w4), .s(w2));   //: @(292, 65) /sz:(51, 50) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>5 Bo0<0 Bo1<0 Bo2<1 ]
  tran g13(.Z(w22), .I(b[11:8]));   //: @(182,13) /sn:0 /R:1 /w:[ 1 6 5 ] /ss:1

endmodule

module main;    //: root_module
wire [15:0] w6;    //: /sn:0 {0}(357,345)(357,401){1}
wire [15:0] w7;    //: /sn:0 {0}(366,213)(366,267){1}
wire w4;    //: /sn:0 {0}(418,345)(418,375){1}
wire [15:0] w0;    //: /sn:0 {0}(457,213)(457,267){1}
wire w1;    //: /sn:0 {0}(497,306)(474,306){1}
wire w2;    //: /sn:0 /dp:1 {0}(334,296)(346,296){1}
wire w5;    //: /sn:0 {0}(442,345)(442,375){1}
//: enddecls

  led g4 (.I(w2));   //: @(327,296) /sn:0 /R:1 /w:[ 0 ] /type:0
  //: frame g8 @(293,183) /sn:0 /wi:249 /ht:262 /tx:""
  //: switch g3 (w1) @(515,306) /sn:0 /R:2 /w:[ 0 ] /st:1
  //: dip g2 (w0) @(457,203) /sn:0 /w:[ 0 ] /st:65535
  //: dip g1 (w7) @(366,203) /sn:0 /w:[ 0 ] /st:65535
  led g6 (.I(w5));   //: @(442,382) /sn:0 /R:2 /w:[ 1 ] /type:0
  led g7 (.I(w4));   //: @(418,382) /sn:0 /R:2 /w:[ 1 ] /type:0
  //: comment g9 /dolink:0 /link:"" @(293,166) /sn:0 /R:2
  //: /line:"Carry Look-Ahead Adder"
  //: /end
  led g5 (.I(w6));   //: @(357,408) /sn:0 /R:2 /w:[ 1 ] /type:3
  CLA16 g0 (.b(w0), .a(w7), .c_in(w1), .c_out(w2), .s(w6), .gg(w5), .pg(w4));   //: @(347, 268) /sz:(126, 76) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<1 Bo0<0 Bo1<0 Bo2<0 ]

endmodule

module CLA(pg, s, b, c_in, a, gg, c_out);
//: interface  /sz:(51, 50) /bd:[ Ti0>a[3:0](14/51) Ti1>b[3:0](33/51) Ri0>c_in(24/50) Bo0<s[3:0](39/51) Bo1<pg(8/51) Bo2<gg(24/51) ]
input [3:0] b;    //: /sn:0 {0}(196,40)(236,40){1}
//: {2}(237,40)(307,40){3}
//: {4}(308,40)(379,40){5}
//: {6}(380,40)(450,40){7}
//: {8}(451,40)(558,40){9}
output pg;    //: /sn:0 {0}(124,259)(424,259)(424,245){1}
output c_out;    //: /sn:0 {0}(125,222)(200,222){1}
input c_in;    //: /sn:0 /dp:1 {0}(468,224)(489,224)(489,109){1}
//: {2}(491,107)(557,107){3}
//: {4}(487,107)(468,107){5}
output [3:0] s;    //: /sn:0 /dp:1 {0}(166,167)(126,167){1}
input [3:0] a;    //: /sn:0 {0}(196,23)(214,23){1}
//: {2}(215,23)(285,23){3}
//: {4}(286,23)(357,23){5}
//: {6}(358,23)(428,23){7}
//: {8}(429,23)(558,23){9}
output gg;    //: /sn:0 {0}(124,274)(442,274)(442,245){1}
wire w16;    //: /sn:0 {0}(297,203)(297,132){1}
wire w13;    //: /sn:0 {0}(451,80)(451,44){1}
wire w25;    //: /sn:0 {0}(308,80)(308,44){1}
wire w22;    //: /sn:0 {0}(424,203)(424,132){1}
wire w36;    //: /sn:0 /dp:1 {0}(172,182)(242,182)(242,132){1}
wire w20;    //: /sn:0 {0}(358,80)(358,27){1}
wire w30;    //: /sn:0 {0}(334,203)(334,107)(325,107){1}
wire w29;    //: /sn:0 {0}(263,203)(263,107)(254,107){1}
wire w12;    //: /sn:0 {0}(281,203)(281,132){1}
wire w18;    //: /sn:0 {0}(456,132)(456,152)(172,152){1}
wire w19;    //: /sn:0 {0}(380,80)(380,44){1}
wire w23;    //: /sn:0 {0}(440,203)(440,132){1}
wire w10;    //: /sn:0 {0}(226,203)(226,132){1}
wire w21;    //: /sn:0 {0}(369,203)(369,132){1}
wire w24;    //: /sn:0 {0}(385,132)(385,162)(172,162){1}
wire w31;    //: /sn:0 {0}(237,80)(237,44){1}
wire w32;    //: /sn:0 {0}(215,80)(215,27){1}
wire w8;    //: /sn:0 {0}(210,203)(210,132){1}
wire w17;    //: /sn:0 {0}(353,203)(353,132){1}
wire w33;    //: /sn:0 {0}(405,203)(405,107)(397,107){1}
wire w14;    //: /sn:0 {0}(429,80)(429,27){1}
wire w15;    //: /sn:0 {0}(172,172)(313,172)(313,132){1}
wire w26;    //: /sn:0 {0}(286,80)(286,27){1}
//: enddecls

  //: output g8 (pg) @(127,259) /sn:0 /R:2 /w:[ 0 ]
  PFA g4 (.a(w32), .b(w31), .c(w29), .s(w36), .g(w10), .p(w8));   //: @(201, 81) /sz:(52, 50) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Bo0<1 Bo1<1 Bo2<1 ]
  PFA g3 (.a(w26), .b(w25), .c(w30), .s(w15), .g(w16), .p(w12));   //: @(272, 81) /sz:(52, 50) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Bo0<1 Bo1<1 Bo2<1 ]
  tran g16(.Z(w32), .I(a[3]));   //: @(215,21) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  //: output g17 (s) @(129,167) /sn:0 /R:2 /w:[ 1 ]
  PFA g2 (.a(w20), .b(w19), .c(w33), .s(w24), .g(w21), .p(w17));   //: @(344, 81) /sz:(52, 50) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Bo0<0 Bo1<1 Bo2<1 ]
  PFA g1 (.a(w14), .b(w13), .c(c_in), .s(w18), .g(w23), .p(w22));   //: @(415, 81) /sz:(52, 50) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>5 Bo0<0 Bo1<1 Bo2<1 ]
  concat g18 (.I0(w18), .I1(w24), .I2(w15), .I3(w36), .Z(s));   //: @(167,167) /sn:0 /R:2 /w:[ 1 1 0 0 0 ] /dr:0
  tran g10(.Z(w19), .I(b[1]));   //: @(380,38) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  //: input g6 (b) @(560,40) /sn:0 /R:2 /w:[ 9 ]
  //: input g7 (c_in) @(559,107) /sn:0 /R:2 /w:[ 3 ]
  tran g9(.Z(w13), .I(b[0]));   //: @(451,38) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  tran g12(.Z(w31), .I(b[3]));   //: @(237,38) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  //: input g5 (a) @(560,23) /sn:0 /R:2 /w:[ 9 ]
  tran g11(.Z(w25), .I(b[2]));   //: @(308,38) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  tran g14(.Z(w20), .I(a[1]));   //: @(358,21) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  //: output g21 (gg) @(127,274) /sn:0 /R:2 /w:[ 0 ]
  //: output g19 (c_out) @(128,222) /sn:0 /R:2 /w:[ 0 ]
  CarryLookaheadLogic g20 (.g0(w23), .p0(w22), .g1(w21), .p1(w17), .g2(w16), .p2(w12), .g3(w10), .p3(w8), .c0(c_in), .c1(w33), .c2(w30), .c3(w29), .c4(c_out), .pg(pg), .gg(gg));   //: @(201, 204) /sz:(266, 40) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>0 Ti3>0 Ti4>0 Ti5>0 Ti6>0 Ti7>0 Ri0>0 To0<0 To1<0 To2<0 Lo0<1 Bo0<1 Bo1<1 ]
  //: joint g0 (c_in) @(489, 107) /w:[ 2 -1 4 1 ]
  tran g15(.Z(w26), .I(a[2]));   //: @(286,21) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  tran g13(.Z(w14), .I(a[0]));   //: @(429,21) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1

endmodule
