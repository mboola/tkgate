//: version "1.8.7"

module main;    //: root_module
wire w4;    //: /sn:0 {0}(358,289)(358,298)(426,298){1}
wire w3;    //: /sn:0 {0}(339,289)(339,333)(456,333)(456,320){1}
wire w0;    //: /sn:0 {0}(452,181)(468,181)(468,278){1}
wire w1;    //: /sn:0 {0}(523,180)(533,180)(533,262)(497,262)(497,298)(485,298){1}
wire w5;    //: /sn:0 {0}(388,181)(400,181)(400,262)(448,262)(448,278){1}
//: enddecls

  led g4 (.I(w4));   //: @(358,282) /sn:0 /w:[ 0 ] /type:0
  //: switch g3 (w1) @(506,180) /sn:0 /w:[ 0 ] /st:0
  //: switch g2 (w0) @(435,181) /sn:0 /w:[ 0 ] /st:0
  //: switch g1 (w5) @(371,181) /sn:0 /w:[ 0 ] /st:0
  led g5 (.I(w3));   //: @(339,282) /sn:0 /w:[ 0 ] /type:0
  FA g0 (.a(w0), .b(w5), .c_in(w1), .c_out(w4), .s(w3));   //: @(427, 279) /sz:(57, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<1 Bo0<1 ]

endmodule

module FA(c_out, s, c_in, b, a);
//: interface  /sz:(57, 40) /bd:[ Ti0>b(21/57) Ti1>a(41/57) Ri0>c_in(19/40) Lo0<c_out(19/40) Bo0<s(29/57) ]
input b;    //: /sn:0 {0}(193,35)(193,98){1}
//: {2}(195,100)(233,100){3}
//: {4}(193,102)(193,162)(300,162){5}
output c_out;    //: /sn:0 /dp:1 {0}(372,145)(398,145){1}
input c_in;    //: /sn:0 /dp:1 {0}(209,35)(209,116){1}
//: {2}(211,118)(282,118)(282,103)(299,103){3}
//: {4}(209,120)(209,144)(300,144){5}
output s;    //: /sn:0 /dp:1 {0}(320,101)(398,101){1}
input a;    //: /sn:0 {0}(177,35)(177,93){1}
//: {2}(179,95)(233,95){3}
//: {4}(177,97)(177,167)(300,167){5}
wire w14;    //: /sn:0 {0}(321,165)(334,165)(334,147)(351,147){1}
wire w11;    //: /sn:0 {0}(321,142)(351,142){1}
wire w2;    //: /sn:0 {0}(254,98)(265,98){1}
//: {2}(269,98)(299,98){3}
//: {4}(267,100)(267,139)(300,139){5}
//: enddecls

  and g8 (.I0(w2), .I1(c_in), .Z(w11));   //: @(311,142) /sn:0 /delay:" 5" /w:[ 5 5 0 ]
  //: output g4 (c_out) @(395,145) /sn:0 /w:[ 1 ]
  //: output g3 (s) @(395,101) /sn:0 /w:[ 1 ]
  //: input g2 (c_in) @(209,33) /sn:0 /R:3 /w:[ 0 ]
  //: input g1 (b) @(193,33) /sn:0 /R:3 /w:[ 0 ]
  //: joint g10 (a) @(177, 95) /w:[ 2 1 -1 4 ]
  xor g6 (.I0(w2), .I1(c_in), .Z(s));   //: @(310,101) /sn:0 /delay:" 6" /w:[ 3 3 0 ]
  and g9 (.I0(b), .I1(a), .Z(w14));   //: @(311,165) /sn:0 /delay:" 5" /w:[ 5 5 0 ]
  or g7 (.I0(w11), .I1(w14), .Z(c_out));   //: @(362,145) /sn:0 /delay:" 5" /w:[ 1 1 0 ]
  //: joint g12 (b) @(193, 100) /w:[ 2 1 -1 4 ]
  xor g5 (.I0(a), .I1(b), .Z(w2));   //: @(244,98) /sn:0 /delay:" 6" /w:[ 3 3 0 ]
  //: joint g11 (w2) @(267, 98) /w:[ 2 -1 1 4 ]
  //: input g0 (a) @(177,33) /sn:0 /R:3 /w:[ 0 ]
  //: joint g13 (c_in) @(209, 118) /w:[ 2 1 -1 4 ]

endmodule
