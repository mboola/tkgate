//: version "1.8.7"

module PFA(p, c, b, g, s, a);
//: interface  /sz:(52, 50) /bd:[ Ti0>a(14/52) Ti1>b(36/52) Ri0>c(26/50) Bo0<s(41/52) Bo1<g(25/52) Bo2<p(9/52) ]
output p;    //: /sn:0 {0}(506,190)(454,190){1}
input b;    //: /sn:0 {0}(265,98)(265,147){1}
//: {2}(267,149)(341,149){3}
//: {4}(265,151)(265,190){5}
//: {6}(267,192)(433,192){7}
//: {8}(265,194)(265,222)(432,222){9}
output s;    //: /sn:0 /dp:1 {0}(453,159)(506,159){1}
input a;    //: /sn:0 {0}(291,98)(291,142){1}
//: {2}(293,144)(341,144){3}
//: {4}(291,146)(291,185){5}
//: {6}(293,187)(433,187){7}
//: {8}(291,189)(291,217)(432,217){9}
output g;    //: /sn:0 {0}(506,220)(453,220){1}
input c;    //: /sn:0 {0}(242,98)(242,161)(432,161){1}
wire w2;    //: /sn:0 {0}(362,147)(393,147)(393,156)(432,156){1}
//: enddecls

  //: output g8 (p) @(503,190) /sn:0 /w:[ 0 ]
  xor g4 (.I0(w2), .I1(c), .Z(s));   //: @(443,159) /sn:0 /delay:" 6" /w:[ 1 1 0 ]
  xor g3 (.I0(a), .I1(b), .Z(w2));   //: @(352,147) /sn:0 /delay:" 6" /w:[ 3 3 0 ]
  //: input g2 (c) @(242,96) /sn:0 /R:3 /w:[ 0 ]
  //: input g1 (b) @(265,96) /sn:0 /R:3 /w:[ 0 ]
  //: joint g10 (a) @(291, 144) /w:[ 2 1 -1 4 ]
  and g6 (.I0(a), .I1(b), .Z(g));   //: @(443,220) /sn:0 /delay:" 5" /w:[ 9 9 1 ]
  //: output g9 (g) @(503,220) /sn:0 /w:[ 0 ]
  //: output g7 (s) @(503,159) /sn:0 /w:[ 1 ]
  //: joint g12 (a) @(291, 187) /w:[ 6 5 -1 8 ]
  //: joint g11 (b) @(265, 192) /w:[ 6 5 -1 8 ]
  or g5 (.I0(a), .I1(b), .Z(p));   //: @(444,190) /sn:0 /delay:" 5" /w:[ 7 7 1 ]
  //: input g0 (a) @(291,96) /sn:0 /R:3 /w:[ 0 ]
  //: joint g13 (b) @(265, 149) /w:[ 2 1 -1 4 ]

endmodule

module main;    //: root_module
wire w6;    //: /sn:0 {0}(345,47)(364,47)(364,160)(413,160)(413,183){1}
wire w4;    //: /sn:0 {0}(424,235)(424,262)(334,262)(334,234){1}
wire w0;    //: /sn:0 {0}(412,47)(435,47)(435,183){1}
wire w1;    //: /sn:0 {0}(493,46)(505,46)(505,165)(475,165)(475,210)(452,210){1}
wire w8;    //: /sn:0 {0}(359,234)(359,270)(440,270)(440,235){1}
wire w5;    //: /sn:0 {0}(408,235)(408,251)(309,251)(309,233){1}
//: enddecls

  led g4 (.I(w5));   //: @(309,226) /sn:0 /w:[ 1 ] /type:0
  //: switch g3 (w1) @(476,46) /sn:0 /w:[ 0 ] /st:0
  //: switch g2 (w0) @(395,47) /sn:0 /w:[ 0 ] /st:0
  //: switch g1 (w6) @(328,47) /sn:0 /w:[ 0 ] /st:0
  led g6 (.I(w8));   //: @(359,227) /sn:0 /w:[ 0 ] /type:0
  led g5 (.I(w4));   //: @(334,227) /sn:0 /w:[ 1 ] /type:0
  PFA g0 (.b(w0), .a(w6), .c(w1), .p(w5), .g(w4), .s(w8));   //: @(399, 184) /sz:(52, 50) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Bo0<0 Bo1<0 Bo2<1 ]

endmodule
