//: version "1.8.7"

module HA(s, b, a, c);
//: interface  /sz:(44, 44) /bd:[ Ti0>b(31/44) Ti1>a(12/44) Lo0<c(20/44) Bo0<s(22/44) ]
input b;    //: /sn:0 /dp:1 {0}(94,103)(125,103)(125,129){1}
//: {2}(127,131)(183,131){3}
//: {4}(125,133)(125,166)(183,166){5}
output s;    //: /sn:0 /dp:1 {0}(204,129)(241,129){1}
input a;    //: /sn:0 /dp:1 {0}(183,161)(137,161)(137,128){1}
//: {2}(139,126)(183,126){3}
//: {4}(137,124)(137,87)(95,87){5}
output c;    //: /sn:0 /dp:1 {0}(204,164)(243,164){1}
//: enddecls

  //: output g4 (s) @(238,129) /sn:0 /w:[ 1 ]
  //: input g3 (b) @(92,103) /sn:0 /w:[ 0 ]
  //: input g2 (a) @(93,87) /sn:0 /w:[ 5 ]
  and g1 (.I0(a), .I1(b), .Z(c));   //: @(194,164) /sn:0 /delay:" 5" /w:[ 0 5 0 ]
  //: joint g6 (b) @(125, 131) /w:[ 2 1 -1 4 ]
  //: joint g7 (a) @(137, 126) /w:[ 2 4 -1 1 ]
  //: output g5 (c) @(240,164) /sn:0 /w:[ 1 ]
  xor g0 (.I0(a), .I1(b), .Z(s));   //: @(194,129) /sn:0 /delay:" 6" /w:[ 3 3 0 ]

endmodule

module main;    //: root_module
wire w4;    //: /sn:0 {0}(358,289)(358,295)(426,295){1}
wire w3;    //: /sn:0 {0}(339,289)(339,333)(449,333)(449,320){1}
wire w0;    //: /sn:0 {0}(452,181)(459,181)(459,273){1}
wire w1;    //: /sn:0 {0}(523,180)(533,180)(533,259)(485,259)(485,295)(473,295){1}
wire w5;    //: /sn:0 {0}(388,181)(395,181)(395,257)(443,257)(443,273){1}
//: enddecls

  led g4 (.I(w4));   //: @(358,282) /sn:0 /w:[ 0 ] /type:0
  //: switch g3 (w1) @(506,180) /sn:0 /w:[ 0 ] /st:1
  //: switch g2 (w0) @(435,181) /sn:0 /w:[ 0 ] /st:1
  //: switch g1 (w5) @(371,181) /sn:0 /w:[ 0 ] /st:1
  led g5 (.I(w3));   //: @(339,282) /sn:0 /w:[ 0 ] /type:0
  FA g0 (.a(w0), .b(w5), .c_in(w1), .c_out(w4), .s(w3));   //: @(427, 274) /sz:(45, 45) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<1 Bo0<1 ]

endmodule

module FA(c_out, s, c_in, b, a);
//: interface  /sz:(57, 40) /bd:[ Ti0>b(21/57) Ti1>a(41/57) Ri0>c_in(19/40) Lo0<c_out(19/40) Bo0<s(29/57) ]
input b;    //: /sn:0 /dp:1 {0}(240,94)(203,94)(203,34){1}
output c_out;    //: /sn:0 /dp:1 {0}(404,147)(427,147){1}
input c_in;    //: /sn:0 {0}(299,37)(299,84)(333,84){1}
output s;    //: /sn:0 {0}(429,93)(379,93){1}
input a;    //: /sn:0 {0}(187,34)(187,113)(240,113){1}
wire w4;    //: /sn:0 /dp:1 {0}(383,149)(261,149)(261,126){1}
wire w0;    //: /sn:0 /dp:1 {0}(383,144)(354,144)(354,116){1}
wire w5;    //: /sn:0 {0}(286,103)(333,103){1}
//: enddecls

  //: output g4 (c_out) @(424,147) /sn:0 /w:[ 1 ]
  //: output g3 (s) @(426,93) /sn:0 /w:[ 0 ]
  //: input g2 (c_in) @(299,35) /sn:0 /R:3 /w:[ 0 ]
  //: input g1 (b) @(203,32) /sn:0 /R:3 /w:[ 1 ]
  or g7 (.I0(w0), .I1(w4), .Z(c_out));   //: @(394,147) /sn:0 /delay:" 5" /w:[ 0 0 0 ]
  HA g14 (.b(b), .a(a), .c(w4), .s(w5));   //: @(241, 81) /sz:(44, 44) /sn:0 /p:[ Li0>0 Li1>1 Bo0<1 Ro0<0 ]
  //: input g0 (a) @(187,32) /sn:0 /R:3 /w:[ 0 ]
  HA g15 (.b(c_in), .a(w5), .c(w0), .s(s));   //: @(334, 71) /sz:(44, 44) /sn:0 /p:[ Li0>1 Li1>1 Bo0<1 Ro0<1 ]

endmodule
