//: version "1.8.7"

module RCA2bits(b, a, s);
//: interface  /sz:(80, 64) /bd:[ Ti0>a[1:0](59/80) Ti1>b[1:0](23/80) Lo0<c(33/64) Bo0<s[1:0](44/80) ]
input [1:0] b;    //: /sn:0 {0}(580,164)(507,164){1}
//: {2}(506,164)(448,164){3}
//: {4}(447,164)(403,164){5}
//: {6}(402,164)(342,164){7}
//: {8}(341,164)(315,164){9}
output [3:0] s;    //: /sn:0 {0}(125,337)(247,337){1}
input [1:0] a;    //: /sn:0 {0}(582,132)(502,132){1}
//: {2}(501,132)(443,132){3}
//: {4}(442,132)(408,132){5}
//: {6}(407,132)(337,132){7}
//: {8}(336,132)(315,132){9}
wire w13;    //: /sn:0 {0}(360,251)(360,234)(390,234)(390,274)(403,274){1}
wire w6;    //: /sn:0 {0}(504,229)(504,322)(253,322){1}
wire w7;    //: /sn:0 {0}(448,168)(448,208){1}
wire w4;    //: /sn:0 {0}(507,168)(507,208){1}
wire w3;    //: /sn:0 {0}(426,299)(426,332)(253,332){1}
wire w0;    //: /sn:0 {0}(416,253)(416,240)(405,240)(405,230){1}
wire w12;    //: /sn:0 /dp:1 {0}(328,272)(312,272)(312,352)(253,352){1}
wire w18;    //: /sn:0 /dp:1 {0}(339,232)(339,251){1}
wire w10;    //: /sn:0 {0}(408,136)(408,209){1}
wire w1;    //: /sn:0 {0}(435,253)(435,240)(445,240)(445,229){1}
wire w8;    //: /sn:0 {0}(443,136)(443,208){1}
wire w2;    //: /sn:0 {0}(342,168)(342,211){1}
wire w11;    //: /sn:0 {0}(403,168)(403,209){1}
wire w15;    //: /sn:0 /dp:1 {0}(351,297)(351,342)(253,342){1}
wire w5;    //: /sn:0 {0}(502,136)(502,208){1}
wire w9;    //: /sn:0 {0}(337,136)(337,211){1}
//: enddecls

  tran g8(.Z(w8), .I(a[1]));   //: @(443,130) /sn:0 /R:1 /w:[ 0 4 3 ] /ss:1
  tran g4(.Z(w4), .I(b[0]));   //: @(507,162) /sn:0 /R:1 /w:[ 0 2 1 ] /ss:1
  tran g16(.Z(w2), .I(b[1]));   //: @(342,162) /sn:0 /R:1 /w:[ 0 8 7 ] /ss:1
  and g3 (.I0(w4), .I1(w5), .Z(w6));   //: @(504,219) /sn:0 /R:3 /delay:" 5" /w:[ 1 1 0 ]
  tran g17(.Z(w9), .I(a[1]));   //: @(337,130) /sn:0 /R:1 /w:[ 0 8 7 ] /ss:1
  //: input g2 (b) @(582,164) /sn:0 /R:2 /w:[ 0 ]
  //: input g1 (a) @(584,132) /sn:0 /R:2 /w:[ 0 ]
  HA g18 (.b(w13), .a(w18), .c(w12), .s(w15));   //: @(329, 252) /sz:(44, 44) /sn:0 /p:[ Ti0>0 Ti1>1 Lo0<0 Bo0<0 ]
  tran g10(.Z(w11), .I(b[1]));   //: @(403,162) /sn:0 /R:1 /w:[ 0 6 5 ] /ss:1
  and g6 (.I0(w7), .I1(w8), .Z(w1));   //: @(445,219) /sn:0 /R:3 /delay:" 5" /w:[ 1 1 1 ]
  and g9 (.I0(w10), .I1(w11), .Z(w0));   //: @(405,220) /sn:0 /R:3 /delay:" 5" /w:[ 1 1 1 ]
  tran g7(.Z(w7), .I(b[0]));   //: @(448,162) /sn:0 /R:1 /w:[ 0 4 3 ] /ss:1
  //: output g12 (s) @(128,337) /sn:0 /R:2 /w:[ 0 ]
  tran g11(.Z(w10), .I(a[0]));   //: @(408,130) /sn:0 /R:1 /w:[ 0 6 5 ] /ss:1
  tran g5(.Z(w5), .I(a[0]));   //: @(502,130) /sn:0 /R:1 /w:[ 0 2 1 ] /ss:1
  and g15 (.I0(w2), .I1(w9), .Z(w18));   //: @(339,222) /sn:0 /R:3 /delay:" 5" /w:[ 1 1 0 ]
  HA g0 (.b(w1), .a(w0), .c(w13), .s(w3));   //: @(404, 254) /sz:(44, 44) /sn:0 /p:[ Ti0>0 Ti1>0 Lo0<1 Bo0<0 ]
  concat g13 (.I0(w6), .I1(w3), .I2(w15), .I3(w12), .Z(s));   //: @(248,337) /sn:0 /R:2 /w:[ 1 1 1 1 1 ] /dr:0

endmodule

module HA(s, b, a, c);
//: interface  /sz:(44, 44) /bd:[ Ti0>a(12/44) Ti1>b(31/44) Lo0<c(20/44) Bo0<s(22/44) ]
input b;    //: /sn:0 /dp:1 {0}(94,103)(125,103)(125,129){1}
//: {2}(127,131)(183,131){3}
//: {4}(125,133)(125,166)(183,166){5}
output s;    //: /sn:0 /dp:1 {0}(204,129)(241,129){1}
input a;    //: /sn:0 /dp:1 {0}(183,161)(137,161)(137,128){1}
//: {2}(139,126)(183,126){3}
//: {4}(137,124)(137,87)(95,87){5}
output c;    //: /sn:0 /dp:1 {0}(204,164)(243,164){1}
//: enddecls

  //: output g4 (s) @(238,129) /sn:0 /w:[ 1 ]
  //: input g3 (b) @(92,103) /sn:0 /w:[ 0 ]
  //: input g2 (a) @(93,87) /sn:0 /w:[ 5 ]
  and g1 (.I0(a), .I1(b), .Z(c));   //: @(194,164) /sn:0 /delay:" 5" /w:[ 0 5 0 ]
  //: joint g6 (b) @(125, 131) /w:[ 2 1 -1 4 ]
  //: joint g7 (a) @(137, 126) /w:[ 2 4 -1 1 ]
  //: output g5 (c) @(240,164) /sn:0 /w:[ 1 ]
  xor g0 (.I0(a), .I1(b), .Z(s));   //: @(194,129) /sn:0 /delay:" 6" /w:[ 3 3 0 ]

endmodule

module main;    //: root_module
wire [3:0] w4;    //: /sn:0 {0}(321,280)(321,322)(414,322)(414,234){1}
wire [1:0] w0;    //: /sn:0 /dp:1 {0}(429,168)(429,121)(460,121)(460,36){1}
wire [1:0] w1;    //: /sn:0 /dp:1 {0}(393,168)(393,123)(359,123)(359,36){1}
//: enddecls

  led g3 (.I(w4));   //: @(321,273) /sn:0 /w:[ 0 ] /type:3
  //: dip g2 (w0) @(460,26) /sn:0 /w:[ 1 ] /st:2
  //: dip g1 (w1) @(359,26) /sn:0 /w:[ 1 ] /st:2
  RCA2bits g0 (.b(w1), .a(w0), .s(w4));   //: @(370, 169) /sz:(80, 64) /sn:0 /p:[ Ti0>0 Ti1>0 Bo0<1 ]

endmodule
