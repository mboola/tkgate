//: version "1.8.7"

module FS(c_in, b, a, c_out, s);
//: interface  /sz:(40, 40) /bd:[ ]
input b;    //: /sn:0 {0}(227,89)(234,89){1}
//: {2}(238,89)(258,89)(258,81)(265,81){3}
//: {4}(236,91)(236,166)(324,166){5}
output c_out;    //: /sn:0 {0}(436,149)(420,149){1}
input c_in;    //: /sn:0 {0}(226,113)(272,113){1}
//: {2}(276,113)(293,113)(293,84)(317,84){3}
//: {4}(274,115)(274,130)(362,130){5}
output s;    //: /sn:0 /dp:1 {0}(338,82)(428,82){1}
input a;    //: /sn:0 {0}(227,76)(239,76){1}
//: {2}(243,76)(265,76){3}
//: {4}(241,78)(241,151)(277,151){5}
wire w7;    //: /sn:0 {0}(383,128)(391,128)(391,146)(399,146){1}
wire w4;    //: /sn:0 {0}(340,117)(354,117)(354,125)(362,125){1}
wire w1;    //: /sn:0 {0}(293,151)(314,151)(314,161)(324,161){1}
wire w2;    //: /sn:0 {0}(286,79)(298,79){1}
//: {2}(302,79)(317,79){3}
//: {4}(300,81)(300,117)(324,117){5}
wire w5;    //: /sn:0 {0}(345,164)(389,164)(389,151)(399,151){1}
//: enddecls

  xor g4 (.I0(w2), .I1(c_in), .Z(s));   //: @(328,82) /sn:0 /delay:" 6" /w:[ 3 3 0 ]
  //: joint g8 (b) @(236, 89) /w:[ 2 -1 1 4 ]
  xor g3 (.I0(a), .I1(b), .Z(w2));   //: @(276,79) /sn:0 /delay:" 6" /w:[ 3 3 0 ]
  //: frame g16 @(184,59) /sn:0 /wi:285 /ht:131 /tx:""
  //: comment g17 /dolink:0 /link:"" @(184,44) /sn:0 /R:2
  //: /line:"Full Substract"
  //: /end
  //: input g2 (c_in) @(224,113) /sn:0 /w:[ 0 ]
  //: input g1 (b) @(225,89) /sn:0 /w:[ 0 ]
  //: joint g10 (w2) @(300, 79) /w:[ 2 -1 1 4 ]
  //: joint g6 (a) @(241, 76) /w:[ 2 -1 1 4 ]
  and g7 (.I0(w1), .I1(b), .Z(w5));   //: @(335,164) /sn:0 /delay:" 5" /w:[ 1 5 0 ]
  not g9 (.I(w2), .Z(w4));   //: @(330,117) /sn:0 /w:[ 5 0 ]
  //: joint g12 (c_in) @(274, 113) /w:[ 2 -1 1 4 ]
  not g5 (.I(a), .Z(w1));   //: @(283,151) /sn:0 /w:[ 5 0 ]
  and g11 (.I0(w4), .I1(c_in), .Z(w7));   //: @(373,128) /sn:0 /delay:" 5" /w:[ 1 5 0 ]
  or g14 (.I0(w7), .I1(w5), .Z(c_out));   //: @(410,149) /sn:0 /delay:" 5" /w:[ 1 1 1 ]
  //: input g0 (a) @(225,76) /sn:0 /w:[ 0 ]
  //: output g15 (c_out) @(433,149) /sn:0 /w:[ 0 ]
  //: output g13 (s) @(425,82) /sn:0 /w:[ 1 ]

endmodule

module CPS4(c_in, a, c_out, s, b);
//: interface  /sz:(40, 40) /bd:[ ]
input [3:0] b;    //: /sn:0 {0}(577,120)(525,120){1}
//: {2}(524,120)(449,120){3}
//: {4}(448,120)(442,120)(442,120)(368,120){5}
//: {6}(367,120)(358,120)(358,120)(275,120){7}
//: {8}(274,120)(248,120){9}
output c_out;    //: /sn:0 /dp:1 {0}(246,174)(219,174){1}
input c_in;    //: /sn:0 {0}(565,179)(540,179){1}
output [3:0] s;    //: /sn:0 /dp:1 {0}(553,235)(593,235){1}
input [3:0] a;    //: /sn:0 {0}(577,100)(507,100){1}
//: {2}(506,100)(484,100)(484,100)(428,100){3}
//: {4}(427,100)(418,100)(418,100)(344,100){5}
//: {6}(343,100)(301,100)(301,100)(258,100){7}
//: {8}(257,100)(243,100){9}
wire w13;    //: /sn:0 {0}(418,176)(376,176){1}
wire w6;    //: /sn:0 {0}(258,104)(258,157){1}
wire w7;    //: /sn:0 {0}(275,124)(275,157){1}
wire w4;    //: /sn:0 {0}(344,104)(344,157){1}
wire w22;    //: /sn:0 /dp:1 {0}(437,203)(437,240)(547,240){1}
wire w3;    //: /sn:0 {0}(449,124)(449,161){1}
wire w0;    //: /sn:0 {0}(507,104)(507,154){1}
wire w12;    //: /sn:0 {0}(498,179)(462,179){1}
wire w23;    //: /sn:0 {0}(353,199)(353,230)(547,230){1}
wire w24;    //: /sn:0 {0}(269,199)(269,220)(547,220){1}
wire w21;    //: /sn:0 /dp:1 {0}(523,198)(523,250)(547,250){1}
wire w1;    //: /sn:0 {0}(525,124)(525,154){1}
wire w14;    //: /sn:0 {0}(333,180)(288,180){1}
wire w2;    //: /sn:0 {0}(428,104)(428,161){1}
wire w5;    //: /sn:0 {0}(368,124)(368,157){1}
//: enddecls

  //: input g8 (c_in) @(567,179) /sn:0 /R:2 /w:[ 0 ]
  //: input g4 (a) @(579,100) /sn:0 /R:2 /w:[ 0 ]
  tran g16(.Z(w6), .I(a[3]));   //: @(258,98) /sn:0 /R:1 /w:[ 0 8 7 ] /ss:1
  FS g3 (.b(w1), .a(w0), .c_in(c_in), .c_out(w12), .s(w21));   //: @(499, 155) /sz:(40, 42) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  //: output g17 (c_out) @(222,174) /sn:0 /R:2 /w:[ 1 ]
  FS g2 (.b(w3), .a(w2), .c_in(w12), .c_out(w13), .s(w22));   //: @(419, 162) /sz:(42, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  //: comment g23 /dolink:0 /link:"" @(530,133) /sn:0
  //: /line:"0T"
  //: /end
  FS g1 (.b(w5), .a(w4), .c_in(w13), .c_out(w14), .s(w23));   //: @(334, 158) /sz:(41, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  //: frame g18 @(174,88) /sn:0 /wi:440 /ht:184 /tx:""
  tran g10(.Z(w0), .I(a[0]));   //: @(507,98) /sn:0 /R:1 /w:[ 0 2 1 ] /ss:1
  concat g6 (.I0(w21), .I1(w22), .I2(w23), .I3(w24), .Z(s));   //: @(552,235) /sn:0 /w:[ 1 1 1 1 0 ] /dr:0
  tran g9(.Z(w1), .I(b[0]));   //: @(525,118) /sn:0 /R:1 /w:[ 0 2 1 ] /ss:1
  //: output g7 (s) @(590,235) /sn:0 /w:[ 1 ]
  //: comment g22 /dolink:0 /link:"" @(499,135) /sn:0
  //: /line:"0T"
  //: /end
  tran g12(.Z(w2), .I(a[1]));   //: @(428,98) /sn:0 /R:1 /w:[ 0 4 3 ] /ss:1
  tran g14(.Z(w4), .I(a[2]));   //: @(344,98) /sn:0 /R:1 /w:[ 0 6 5 ] /ss:1
  tran g11(.Z(w3), .I(b[1]));   //: @(449,118) /sn:0 /R:1 /w:[ 0 4 3 ] /ss:1
  //: input g5 (b) @(579,120) /sn:0 /R:2 /w:[ 0 ]
  //: comment g19 /dolink:0 /link:"" @(175,70) /sn:0 /R:2
  //: /line:"Carry Propagate Substract 4bits"
  //: /end
  //: comment g21 /dolink:0 /link:"" @(561,163) /sn:0
  //: /line:"0T"
  //: /end
  tran g15(.Z(w7), .I(b[3]));   //: @(275,118) /sn:0 /R:1 /w:[ 0 8 7 ] /ss:1
  FS g0 (.b(w7), .a(w6), .c_in(w14), .c_out(c_out), .s(w24));   //: @(247, 158) /sz:(40, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  tran g13(.Z(w5), .I(b[2]));   //: @(368,118) /sn:0 /R:1 /w:[ 0 6 5 ] /ss:1

endmodule

module CPS16(c_in, s, b, c_out, a);
//: interface  /sz:(101, 91) /bd:[ ]
input [15:0] b;    //: /sn:0 {0}(115,123)(207,123){1}
//: {2}(208,123)(350,123){3}
//: {4}(351,123)(478,123){5}
//: {6}(479,123)(604,123){7}
//: {8}(605,123)(634,123){9}
output c_out;    //: /sn:0 {0}(124,227)(154,227){1}
input c_in;    //: /sn:0 {0}(666,219)(619,219){1}
output [15:0] s;    //: /sn:0 {0}(666,317)(701,317){1}
input [15:0] a;    //: /sn:0 {0}(116,149)(175,149){1}
//: {2}(176,149)(316,149){3}
//: {4}(317,149)(436,149){5}
//: {6}(437,149)(572,149){7}
//: {8}(573,149)(625,149){9}
wire [3:0] w16;    //: /sn:0 {0}(605,127)(605,182){1}
wire [3:0] w13;    //: /sn:0 {0}(485,246)(485,322)(660,322){1}
wire [3:0] w6;    //: /sn:0 {0}(351,127)(351,191){1}
wire [3:0] w4;    //: /sn:0 {0}(317,153)(317,191){1}
wire [3:0] w3;    //: /sn:0 /dp:1 {0}(176,189)(176,153){1}
wire [3:0] w0;    //: /sn:0 /dp:1 {0}(208,189)(208,127){1}
wire [3:0] w12;    //: /sn:0 {0}(607,242)(607,302)(660,302){1}
wire w19;    //: /sn:0 {0}(555,220)(502,220){1}
wire [3:0] w10;    //: /sn:0 {0}(437,153)(437,181){1}
wire [3:0] w1;    //: /sn:0 {0}(192,253)(192,332)(660,332){1}
wire [3:0] w8;    //: /sn:0 /dp:1 {0}(346,244)(346,312)(660,312){1}
wire w14;    //: /sn:0 {0}(420,220)(365,220){1}
wire [3:0] w11;    //: /sn:0 {0}(479,127)(479,181){1}
wire [3:0] w15;    //: /sn:0 {0}(573,153)(573,182){1}
wire w9;    //: /sn:0 {0}(302,216)(225,216){1}
//: enddecls

  //: input g4 (c_in) @(668,219) /sn:0 /R:2 /w:[ 0 ]
  //: output g8 (s) @(698,317) /sn:0 /w:[ 1 ]
  tran g16(.Z(w0), .I(b[15:12]));   //: @(208,121) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  CPS4 g3 (.b(w16), .a(w15), .c_in(c_in), .c_out(w19), .s(w12));   //: @(556, 183) /sz:(62, 58) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  tran g17(.Z(w3), .I(a[15:12]));   //: @(176,147) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  CPS4 g2 (.b(w11), .a(w10), .c_in(w19), .c_out(w14), .s(w13));   //: @(421, 182) /sz:(80, 63) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  CPS4 g1 (.b(w6), .a(w4), .c_in(w14), .c_out(w9), .s(w8));   //: @(303, 192) /sz:(61, 51) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  //: frame g18 @(89,104) /sn:0 /wi:626 /ht:246 /tx:""
  tran g10(.Z(w16), .I(b[3:0]));   //: @(605,121) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  //: input g6 (b) @(113,123) /sn:0 /w:[ 0 ]
  concat g7 (.I0(w12), .I1(w8), .I2(w13), .I3(w1), .Z(s));   //: @(665,317) /sn:0 /w:[ 1 1 1 1 0 ] /dr:1
  //: output g9 (c_out) @(127,227) /sn:0 /R:2 /w:[ 0 ]
  tran g12(.Z(w11), .I(b[7:4]));   //: @(479,121) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  tran g14(.Z(w4), .I(a[11:8]));   //: @(317,147) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  tran g11(.Z(w15), .I(a[3:0]));   //: @(573,147) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  //: input g5 (a) @(114,149) /sn:0 /w:[ 0 ]
  //: comment g19 /dolink:0 /link:"" @(90,83) /sn:0 /R:2
  //: /line:"Carry Propagate Substract"
  //: /end
  tran g15(.Z(w10), .I(a[7:4]));   //: @(437,147) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  CPS4 g0 (.b(w0), .a(w3), .c_in(w9), .c_out(c_out), .s(w1));   //: @(155, 190) /sz:(69, 62) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<1 Bo0<0 ]
  tran g13(.Z(w6), .I(b[11:8]));   //: @(351,121) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1

endmodule

module main;    //: root_module
wire [15:0] w4;    //: /sn:0 {0}(213,223)(213,173){1}
wire [15:0] w0;    //: /sn:0 /dp:1 {0}(176,48)(176,80){1}
wire w3;    //: /sn:0 {0}(120,129)(156,129){1}
wire [15:0] w2;    //: /sn:0 /dp:1 {0}(235,22)(235,80){1}
wire w5;    //: /sn:0 {0}(301,128)(259,128){1}
//: enddecls

  //: dip g4 (w0) @(176,38) /sn:0 /w:[ 0 ] /st:10
  led g3 (.I(w4));   //: @(213,230) /sn:0 /R:2 /w:[ 0 ] /type:3
  led g2 (.I(w3));   //: @(113,129) /sn:0 /R:1 /w:[ 0 ] /type:0
  //: switch g1 (w5) @(319,128) /sn:0 /R:2 /w:[ 0 ] /st:0
  //: frame g6 @(94,-4) /sn:0 /wi:251 /ht:270 /tx:""
  //: comment g7 /dolink:0 /link:"" @(95,-18) /sn:0 /R:2
  //: /line:"Carry Propagate Substract"
  //: /end
  //: dip g5 (w2) @(235,12) /sn:0 /w:[ 0 ] /st:2
  CPS16 g0 (.a(w0), .b(w2), .c_in(w5), .c_out(w3), .s(w4));   //: @(157, 81) /sz:(101, 91) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<1 Bo0<1 ]

endmodule
