//: version "1.8.7"

module CPA(c_out, s, c_in, b, a);
//: interface  /sz:(90, 79) /bd:[ Ti0>a[3:0](24/90) Ti1>b[3:0](67/90) Ri0>c_in(40/79) Lo0<c_out(41/79) Bo0<s[3:0](46/90) ]
input [3:0] b;    //: /sn:0 {0}(548,173)(428,173){1}
//: {2}(427,173)(342,173){3}
//: {4}(341,173)(257,173){5}
//: {6}(256,173)(170,173){7}
//: {8}(169,173)(148,173){9}
output c_out;    //: /sn:0 {0}(53,269)(148,269){1}
input c_in;    //: /sn:0 {0}(549,214)(483,214)(483,269)(465,269){1}
output [3:0] s;    //: /sn:0 /dp:1 {0}(102,326)(83,326)(83,286)(53,286){1}
input [3:0] a;    //: /sn:0 {0}(548,191)(448,191){1}
//: {2}(447,191)(362,191){3}
//: {4}(361,191)(277,191){5}
//: {6}(276,191)(190,191){7}
//: {8}(189,191)(148,191){9}
wire w16;    //: /sn:0 {0}(170,249)(170,177){1}
wire w6;    //: /sn:0 {0}(342,249)(342,177){1}
wire w22;    //: /sn:0 /dp:1 {0}(108,341)(178,341)(178,291){1}
wire w3;    //: /sn:0 {0}(406,269)(379,269){1}
wire w0;    //: /sn:0 {0}(448,249)(448,195){1}
wire w20;    //: /sn:0 /dp:1 {0}(108,311)(436,311)(436,291){1}
wire w18;    //: /sn:0 /dp:1 {0}(108,321)(350,321)(350,291){1}
wire w12;    //: /sn:0 {0}(294,269)(320,269){1}
wire w10;    //: /sn:0 {0}(277,249)(277,195){1}
wire w1;    //: /sn:0 {0}(428,249)(428,177){1}
wire w8;    //: /sn:0 /dp:1 {0}(108,331)(265,331)(265,291){1}
wire w17;    //: /sn:0 {0}(207,269)(235,269){1}
wire w11;    //: /sn:0 {0}(257,249)(257,177){1}
wire w15;    //: /sn:0 {0}(190,249)(190,195){1}
wire w5;    //: /sn:0 {0}(362,249)(362,195){1}
//: enddecls

  FA g8 (.b(w16), .a(w15), .c_in(w17), .c_out(c_out), .s(w22));   //: @(149, 250) /sz:(57, 40) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>0 Lo0<1 Bo0<1 ]
  //: output g4 (c_out) @(56,269) /sn:0 /R:2 /w:[ 0 ]
  tran g16(.Z(w11), .I(b[2]));   //: @(257,171) /sn:0 /R:1 /w:[ 1 6 5 ] /ss:1
  //: output g3 (s) @(56,286) /sn:0 /R:2 /w:[ 1 ]
  tran g17(.Z(w16), .I(b[3]));   //: @(170,171) /sn:0 /R:1 /w:[ 1 8 7 ] /ss:1
  //: input g2 (c_in) @(551,214) /sn:0 /R:2 /w:[ 0 ]
  //: input g1 (b) @(550,173) /sn:0 /R:2 /w:[ 0 ]
  tran g10(.Z(w0), .I(a[0]));   //: @(448,189) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:1
  FA g6 (.b(w6), .a(w5), .c_in(w3), .c_out(w12), .s(w18));   //: @(321, 250) /sz:(57, 40) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<1 Bo0<1 ]
  concat g9 (.I0(w20), .I1(w18), .I2(w8), .I3(w22), .Z(s));   //: @(103,326) /sn:0 /R:2 /w:[ 0 0 0 0 0 ] /dr:0
  FA g7 (.b(w11), .a(w10), .c_in(w12), .c_out(w17), .s(w8));   //: @(236, 250) /sz:(57, 40) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>0 Lo0<1 Bo0<1 ]
  tran g12(.Z(w10), .I(a[2]));   //: @(277,189) /sn:0 /R:1 /w:[ 1 6 5 ] /ss:1
  tran g14(.Z(w1), .I(b[0]));   //: @(428,171) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:1
  tran g11(.Z(w5), .I(a[1]));   //: @(362,189) /sn:0 /R:1 /w:[ 1 4 3 ] /ss:1
  FA g5 (.b(w1), .a(w0), .c_in(c_in), .c_out(w3), .s(w20));   //: @(407, 250) /sz:(57, 40) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<0 Bo0<1 ]
  tran g15(.Z(w6), .I(b[1]));   //: @(342,171) /sn:0 /R:1 /w:[ 1 4 3 ] /ss:1
  //: input g0 (a) @(550,191) /sn:0 /R:2 /w:[ 0 ]
  tran g13(.Z(w15), .I(a[3]));   //: @(190,189) /sn:0 /R:1 /w:[ 1 8 7 ] /ss:1

endmodule

module FA(c_out, s, c_in, b, a);
//: interface  /sz:(85, 65) /bd:[ Ti0>a(19/85) Ti1>b(68/85) Ri0>c_in(33/65) Lo0<c_out(32/65) Bo0<s(43/85) ]
input b;    //: /sn:0 {0}(188,79)(188,149){1}
//: {2}(190,151)(247,151){3}
//: {4}(188,153)(188,225){5}
//: {6}(190,227)(247,227){7}
//: {8}(188,229)(188,261)(247,261){9}
output c_out;    //: /sn:0 /dp:1 {0}(393,213)(423,213){1}
input c_in;    //: /sn:0 {0}(206,79)(206,164){1}
//: {2}(208,166)(295,166)(295,154)(314,154){3}
//: {4}(206,168)(206,190){5}
//: {6}(208,192)(247,192){7}
//: {8}(206,194)(206,256)(247,256){9}
output s;    //: /sn:0 /dp:1 {0}(335,152)(423,152){1}
input a;    //: /sn:0 {0}(171,79)(171,144){1}
//: {2}(173,146)(247,146){3}
//: {4}(171,148)(171,185){5}
//: {6}(173,187)(247,187){7}
//: {8}(171,189)(171,222)(247,222){9}
wire w7;    //: /sn:0 {0}(268,259)(352,259)(352,215)(372,215){1}
wire w4;    //: /sn:0 {0}(268,190)(296,190)(296,207)(315,207){1}
wire w0;    //: /sn:0 /dp:1 {0}(314,149)(268,149){1}
wire w8;    //: /sn:0 {0}(336,210)(372,210){1}
wire w5;    //: /sn:0 {0}(268,225)(296,225)(296,212)(315,212){1}
//: enddecls

  xor g8 (.I0(w0), .I1(c_in), .Z(s));   //: @(325,152) /sn:0 /delay:" 6" /w:[ 0 3 0 ]
  //: output g4 (c_out) @(420,213) /sn:0 /w:[ 1 ]
  or g16 (.I0(w4), .I1(w5), .Z(w8));   //: @(326,210) /sn:0 /delay:" 5" /w:[ 1 1 0 ]
  //: output g3 (s) @(420,152) /sn:0 /w:[ 1 ]
  or g17 (.I0(w8), .I1(w7), .Z(c_out));   //: @(383,213) /sn:0 /delay:" 5" /w:[ 1 1 0 ]
  //: input g2 (c_in) @(206,77) /sn:0 /R:3 /w:[ 0 ]
  //: input g1 (b) @(188,77) /sn:0 /R:3 /w:[ 0 ]
  and g10 (.I0(a), .I1(c_in), .Z(w4));   //: @(258,190) /sn:0 /delay:" 5" /w:[ 7 7 0 ]
  xor g6 (.I0(a), .I1(b), .Z(w0));   //: @(258,149) /sn:0 /delay:" 6" /w:[ 3 3 1 ]
  //: joint g7 (b) @(188, 151) /w:[ 2 1 -1 4 ]
  //: joint g9 (a) @(171, 146) /w:[ 2 1 -1 4 ]
  //: joint g12 (c_in) @(206, 192) /w:[ 6 5 -1 8 ]
  //: joint g14 (b) @(188, 227) /w:[ 6 5 -1 8 ]
  //: joint g11 (a) @(171, 187) /w:[ 6 5 -1 8 ]
  //: joint g5 (c_in) @(206, 166) /w:[ 2 1 -1 4 ]
  and g15 (.I0(c_in), .I1(b), .Z(w7));   //: @(258,259) /sn:0 /delay:" 5" /w:[ 9 9 0 ]
  //: input g0 (a) @(171,77) /sn:0 /R:3 /w:[ 0 ]
  and g13 (.I0(a), .I1(b), .Z(w5));   //: @(258,225) /sn:0 /delay:" 5" /w:[ 9 7 0 ]

endmodule

module main;    //: root_module
wire [4:0] w6;    //: /sn:0 {0}(435,243)(435,326)(386,326){1}
wire w4;    //: /sn:0 {0}(260,255)(237,255)(237,321)(380,321){1}
wire [3:0] w0;    //: /sn:0 /dp:1 {0}(285,213)(285,171)(187,171)(187,86){1}
wire w1;    //: /sn:0 {0}(363,75)(387,75)(387,254)(352,254){1}
wire [3:0] w2;    //: /sn:0 {0}(307,294)(307,331)(380,331){1}
wire [3:0] w5;    //: /sn:0 {0}(276,86)(276,139)(328,139)(328,213){1}
//: enddecls

  concat g4 (.I0(w2), .I1(w4), .Z(w6));   //: @(385,326) /sn:0 /w:[ 1 1 1 ] /dr:0
  //: switch g3 (w1) @(346,75) /sn:0 /w:[ 0 ] /st:0
  //: dip g2 (w0) @(187,76) /sn:0 /w:[ 1 ] /st:15
  //: dip g1 (w5) @(276,76) /sn:0 /w:[ 0 ] /st:15
  led g5 (.I(w6));   //: @(435,236) /sn:0 /w:[ 0 ] /type:3
  CPA g0 (.b(w5), .a(w0), .c_in(w1), .c_out(w4), .s(w2));   //: @(261, 214) /sz:(90, 79) /sn:0 /p:[ Ti0>1 Ti1>0 Ri0>1 Lo0<0 Bo0<0 ]

endmodule
