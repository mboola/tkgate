//: version "1.8.7"

module RCA4bits(s, b, a);
//: interface  /sz:(77, 73) /bd:[ Ti0>b[3:0](57/77) Ti1>a[3:0](22/77) Bo0<s[6:0](38/77) ]
input [3:0] b;    //: /sn:0 {0}(798,-233)(798,-216){1}
//: {2}(798,-215)(798,-84){3}
//: {4}(798,-83)(798,128){5}
//: {6}(798,129)(798,301){7}
//: {8}(798,302)(798,351){9}
output [7:0] s;    //: /sn:0 {0}(-105,522)(-12,522){1}
input [3:0] a;    //: /sn:0 {0}(738,-343)(702,-343){1}
//: {2}(701,-343)(668,-343){3}
//: {4}(667,-343)(630,-343){5}
//: {6}(629,-343)(595,-343){7}
//: {8}(594,-343)(575,-343){9}
wire w13;    //: /sn:0 {0}(785,129)(390,129){1}
//: {2}(386,129)(309,129){3}
//: {4}(305,129)(237,129){5}
//: {6}(233,129)(161,129)(161,193){7}
//: {8}(235,131)(235,193){9}
//: {10}(307,131)(307,193){11}
//: {12}(388,131)(388,192){13}
wire w58;    //: /sn:0 {0}(222,100)(222,235){1}
wire w7;    //: /sn:0 /dp:1 {0}(172,369)(172,331)(630,331)(630,162){1}
//: {2}(630,158)(630,-42){3}
//: {4}(630,-46)(630,-186){5}
//: {6}(630,-190)(630,-339){7}
//: {8}(628,-188)(368,-188)(368,-145){9}
//: {10}(628,-44)(306,-44)(306,-6){11}
//: {12}(628,160)(240,160)(240,193){13}
wire w34;    //: /sn:0 {0}(211,432)(183,432){1}
wire w59;    //: /sn:0 {0}(288,-124)(288,53){1}
wire w72;    //: /sn:0 {0}(163,214)(163,235){1}
wire w0;    //: /sn:0 {0}(785,-215)(513,-215){1}
//: {2}(509,-215)(440,-215){3}
//: {4}(436,-215)(365,-215){5}
//: {6}(361,-215)(286,-215)(286,-145){7}
//: {8}(363,-213)(363,-145){9}
//: {10}(438,-213)(438,-145){11}
//: {12}(511,-213)(511,-145){13}
wire w3;    //: /sn:0 {0}(440,53)(440,-124){1}
wire w22;    //: /sn:0 {0}(459,15)(459,53){1}
wire w36;    //: /sn:0 {0}(394,74)(427,74){1}
wire w20;    //: /sn:0 {0}(450,99)(450,497)(-6,497){1}
wire w30;    //: /sn:0 {0}(287,432)(257,432){1}
wire w29;    //: /sn:0 /dp:1 {0}(246,369)(246,345)(668,345)(668,175){1}
//: {2}(668,171)(668,-27){3}
//: {4}(668,-31)(668,-171){5}
//: {6}(668,-175)(668,-339){7}
//: {8}(666,-173)(443,-173)(443,-145){9}
//: {10}(666,-29)(383,-29)(383,-7){11}
//: {12}(666,173)(312,173)(312,193){13}
wire w37;    //: /sn:0 {0}(137,432)(110,432){1}
wire w42;    //: /sn:0 {0}(371,99)(371,235){1}
wire w66;    //: /sn:0 {0}(390,213)(390,235){1}
wire w63;    //: /sn:0 {0}(303,15)(303,53){1}
wire w54;    //: /sn:0 {0}(154,281)(154,411){1}
wire w70;    //: /sn:0 {0}(237,214)(237,235){1}
wire w1;    //: /sn:0 {0}(702,-339)(702,-153){1}
//: {2}(700,-151)(516,-151)(516,-145){3}
//: {4}(702,-149)(702,-18){5}
//: {6}(700,-16)(462,-16)(462,-6){7}
//: {8}(702,-14)(702,184){9}
//: {10}(700,186)(393,186)(393,192){11}
//: {12}(702,188)(702,359)(322,359)(322,369){13}
wire w31;    //: /sn:0 {0}(310,457)(310,517)(-6,517){1}
wire w68;    //: /sn:0 {0}(309,214)(309,235){1}
wire w53;    //: /sn:0 {0}(131,256)(81,256)(81,411){1}
wire w46;    //: /sn:0 {0}(300,281)(300,411){1}
wire w8;    //: /sn:0 /dp:1 {0}(99,370)(99,317)(595,317)(595,148){1}
//: {2}(595,144)(595,-59){3}
//: {4}(595,-63)(595,-201){5}
//: {6}(595,-205)(595,-339){7}
//: {8}(593,-203)(291,-203)(291,-145){9}
//: {10}(593,-61)(215,-61)(215,-4){11}
//: {12}(593,146)(166,146)(166,193){13}
wire w52;    //: /sn:0 {0}(294,99)(294,235){1}
wire w44;    //: /sn:0 {0}(323,256)(358,256){1}
wire w28;    //: /sn:0 {0}(381,281)(381,507)(-6,507){1}
wire w35;    //: /sn:0 {0}(234,457)(234,527)(-6,527){1}
wire w80;    //: /sn:0 {0}(96,391)(96,411){1}
wire w45;    //: /sn:0 {0}(277,256)(251,256){1}
wire w49;    //: /sn:0 {0}(228,281)(228,411){1}
wire w2;    //: /sn:0 {0}(513,-124)(513,487)(-6,487){1}
wire w11;    //: /sn:0 {0}(785,-83)(459,-83){1}
//: {2}(455,-83)(380,-83){3}
//: {4}(376,-83)(303,-83){5}
//: {6}(299,-83)(210,-83)(210,-4){7}
//: {8}(301,-81)(301,-6){9}
//: {10}(378,-81)(378,-7){11}
//: {12}(457,-81)(457,-6){13}
wire w48;    //: /sn:0 {0}(205,256)(177,256){1}
wire w41;    //: /sn:0 {0}(365,-124)(365,53){1}
wire w74;    //: /sn:0 {0}(319,390)(319,411){1}
wire w78;    //: /sn:0 {0}(169,390)(169,411){1}
wire w47;    //: /sn:0 {0}(271,74)(256,74)(256,44)(231,44)(231,54){1}
wire w15;    //: /sn:0 {0}(785,302)(319,302){1}
//: {2}(315,302)(243,302){3}
//: {4}(239,302)(169,302){5}
//: {6}(165,302)(94,302)(94,370){7}
//: {8}(167,304)(167,369){9}
//: {10}(241,304)(241,369){11}
//: {12}(317,304)(317,369){13}
wire w38;    //: /sn:0 {0}(160,457)(160,537)(-6,537){1}
wire w61;    //: /sn:0 {0}(212,17)(212,54){1}
wire w43;    //: /sn:0 {0}(87,457)(87,547)(-6,547){1}
wire w64;    //: /sn:0 {0}(380,14)(380,53){1}
wire w9;    //: /sn:0 {0}(-6,557)(47,557)(47,432)(64,432){1}
wire w76;    //: /sn:0 {0}(243,390)(243,411){1}
wire w40;    //: /sn:0 {0}(317,74)(348,74){1}
wire w57;    //: /sn:0 {0}(199,75)(148,75)(148,235){1}
//: enddecls

  concat g4 (.I0(w2), .I1(w20), .I2(w28), .I3(w31), .I4(w35), .I5(w38), .I6(w43), .I7(w9), .Z(s));   //: @(-11,522) /sn:0 /R:2 /w:[ 1 1 1 1 1 1 1 0 1 ] /dr:0
  tran g8(.Z(w29), .I(a[1]));   //: @(668,-345) /sn:0 /R:1 /w:[ 7 4 3 ] /ss:1
  //: joint g44 (w13) @(307, 129) /w:[ 3 -1 4 10 ]
  and g3 (.I0(w1), .I1(w0), .Z(w2));   //: @(513,-134) /sn:0 /R:3 /delay:" 5" /w:[ 3 13 0 ]
  HA g16 (.b(w74), .a(w46), .c(w30), .s(w31));   //: @(288, 412) /sz:(44, 44) /sn:0 /p:[ Ti0>1 Ti1>1 Lo0<0 Bo0<0 ]
  //: joint g47 (w11) @(378, -83) /w:[ 3 -1 4 10 ]
  FA g17 (.b(w49), .a(w76), .c_in(w30), .c_out(w34), .s(w35));   //: @(212, 412) /sz:(44, 44) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  HA g26 (.b(w47), .a(w61), .c(w57), .s(w58));   //: @(200, 55) /sz:(44, 44) /sn:0 /p:[ Ti0>1 Ti1>1 Lo0<0 Bo0<0 ]
  //: output g2 (s) @(-102,522) /sn:0 /R:2 /w:[ 0 ]
  FA g23 (.b(w58), .a(w70), .c_in(w45), .c_out(w48), .s(w49));   //: @(206, 236) /sz:(44, 44) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  and g30 (.I0(w7), .I1(w11), .Z(w63));   //: @(303,5) /sn:0 /R:3 /delay:" 5" /w:[ 11 9 0 ]
  //: input g1 (b) @(798,-235) /sn:0 /R:3 /w:[ 0 ]
  FA g24 (.b(w57), .a(w72), .c_in(w48), .c_out(w53), .s(w54));   //: @(132, 236) /sz:(44, 44) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  and g39 (.I0(w8), .I1(w15), .Z(w80));   //: @(96,381) /sn:0 /R:3 /delay:" 5" /w:[ 0 7 0 ]
  and g29 (.I0(w8), .I1(w11), .Z(w61));   //: @(212,7) /sn:0 /R:3 /delay:" 5" /w:[ 11 7 0 ]
  //: joint g60 (w1) @(702, -151) /w:[ -1 1 2 4 ]
  //: joint g51 (w0) @(363, -215) /w:[ 5 -1 6 8 ]
  FA g18 (.b(w54), .a(w78), .c_in(w34), .c_out(w37), .s(w38));   //: @(138, 412) /sz:(44, 44) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  tran g10(.Z(w7), .I(a[2]));   //: @(630,-345) /sn:0 /R:1 /w:[ 7 6 5 ] /ss:1
  FA g25 (.b(w59), .a(w63), .c_in(w40), .c_out(w47), .s(w52));   //: @(272, 54) /sz:(44, 44) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<0 Bo0<0 ]
  //: joint g49 (w0) @(511, -215) /w:[ 1 -1 2 12 ]
  tran g6(.Z(w1), .I(a[0]));   //: @(702,-345) /sn:0 /R:1 /w:[ 0 2 1 ] /ss:1
  //: joint g50 (w0) @(438, -215) /w:[ 3 -1 4 10 ]
  tran g7(.Z(w11), .I(b[1]));   //: @(796,-83) /sn:0 /R:2 /w:[ 0 4 3 ] /ss:0
  tran g9(.Z(w13), .I(b[2]));   //: @(796,129) /sn:0 /R:2 /w:[ 0 6 5 ] /ss:0
  and g35 (.I0(w8), .I1(w13), .Z(w72));   //: @(163,204) /sn:0 /R:3 /delay:" 5" /w:[ 13 7 0 ]
  //: joint g56 (w8) @(595, 146) /w:[ -1 2 12 1 ]
  //: joint g58 (w29) @(668, 173) /w:[ -1 2 12 1 ]
  FA g22 (.b(w52), .a(w68), .c_in(w44), .c_out(w45), .s(w46));   //: @(278, 236) /sz:(44, 44) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<0 Bo0<0 ]
  and g31 (.I0(w29), .I1(w11), .Z(w64));   //: @(380,4) /sn:0 /R:3 /delay:" 5" /w:[ 11 11 0 ]
  //: joint g59 (w1) @(702, 186) /w:[ -1 9 10 12 ]
  and g33 (.I0(w29), .I1(w13), .Z(w68));   //: @(309,204) /sn:0 /R:3 /delay:" 5" /w:[ 13 11 0 ]
  and g36 (.I0(w1), .I1(w15), .Z(w74));   //: @(319,380) /sn:0 /R:3 /delay:" 5" /w:[ 13 13 0 ]
  //: joint g41 (w15) @(241, 302) /w:[ 3 -1 4 10 ]
  //: joint g45 (w13) @(235, 129) /w:[ 5 -1 6 8 ]
  //: joint g54 (w29) @(668, -29) /w:[ -1 4 10 3 ]
  //: joint g40 (w15) @(317, 302) /w:[ 1 -1 2 12 ]
  //: joint g42 (w15) @(167, 302) /w:[ 5 -1 6 8 ]
  //: joint g52 (w8) @(595, -61) /w:[ -1 4 10 3 ]
  tran g12(.Z(w8), .I(a[3]));   //: @(595,-345) /sn:0 /R:1 /w:[ 7 8 7 ] /ss:1
  and g28 (.I0(w8), .I1(w0), .Z(w59));   //: @(288,-134) /sn:0 /R:3 /delay:" 5" /w:[ 9 7 0 ]
  and g34 (.I0(w7), .I1(w13), .Z(w70));   //: @(237,204) /sn:0 /R:3 /delay:" 5" /w:[ 13 9 0 ]
  //: joint g46 (w11) @(457, -83) /w:[ 1 -1 2 12 ]
  //: joint g57 (w7) @(630, 160) /w:[ -1 2 12 1 ]
  tran g5(.Z(w0), .I(b[0]));   //: @(796,-215) /sn:0 /R:2 /w:[ 0 2 1 ] /ss:0
  tran g11(.Z(w15), .I(b[3]));   //: @(796,302) /sn:0 /R:2 /w:[ 0 8 7 ] /ss:0
  and g14 (.I0(w1), .I1(w11), .Z(w22));   //: @(459,5) /sn:0 /R:3 /delay:" 5" /w:[ 7 13 0 ]
  FA g19 (.b(w53), .a(w80), .c_in(w37), .c_out(w9), .s(w43));   //: @(65, 412) /sz:(44, 44) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<1 Bo0<0 ]
  FA g21 (.b(w41), .a(w64), .c_in(w36), .c_out(w40), .s(w42));   //: @(349, 54) /sz:(44, 44) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  //: joint g61 (w29) @(668, -173) /w:[ -1 6 8 5 ]
  and g20 (.I0(w29), .I1(w0), .Z(w3));   //: @(440,-134) /sn:0 /R:3 /delay:" 5" /w:[ 9 11 1 ]
  and g32 (.I0(w1), .I1(w13), .Z(w66));   //: @(390,203) /sn:0 /R:3 /delay:" 5" /w:[ 11 13 0 ]
  //: joint g63 (w8) @(595, -203) /w:[ -1 6 8 5 ]
  //: input g0 (a) @(740,-343) /sn:0 /R:2 /w:[ 0 ]
  HA g15 (.b(w66), .a(w42), .c(w44), .s(w28));   //: @(359, 236) /sz:(44, 44) /sn:0 /p:[ Ti0>1 Ti1>1 Lo0<1 Bo0<0 ]
  and g38 (.I0(w7), .I1(w15), .Z(w78));   //: @(169,380) /sn:0 /R:3 /delay:" 5" /w:[ 0 9 0 ]
  //: joint g43 (w13) @(388, 129) /w:[ 1 -1 2 12 ]
  and g27 (.I0(w7), .I1(w0), .Z(w41));   //: @(365,-134) /sn:0 /R:3 /delay:" 5" /w:[ 9 9 0 ]
  //: joint g48 (w11) @(301, -83) /w:[ 5 -1 6 8 ]
  and g37 (.I0(w29), .I1(w15), .Z(w76));   //: @(243,380) /sn:0 /R:3 /delay:" 5" /w:[ 0 11 0 ]
  //: joint g62 (w7) @(630, -188) /w:[ -1 6 8 5 ]
  //: joint g55 (w1) @(702, -16) /w:[ -1 5 6 8 ]
  HA g13 (.b(w22), .a(w3), .c(w36), .s(w20));   //: @(428, 54) /sz:(44, 44) /sn:0 /p:[ Ti0>1 Ti1>0 Lo0<1 Bo0<0 ]
  //: joint g53 (w7) @(630, -44) /w:[ -1 4 10 3 ]

endmodule

module HA(s, b, a, c);
//: interface  /sz:(44, 44) /bd:[ Ti0>a(12/44) Ti1>b(31/44) Ti2>b(31/44) Ti3>a(12/44) Lo0<c(20/44) Lo1<c(20/44) Bo0<s(22/44) Bo1<s(22/44) ]
input b;    //: /sn:0 /dp:1 {0}(94,103)(125,103)(125,129){1}
//: {2}(127,131)(183,131){3}
//: {4}(125,133)(125,166)(183,166){5}
output s;    //: /sn:0 /dp:1 {0}(204,129)(241,129){1}
input a;    //: /sn:0 /dp:1 {0}(183,161)(137,161)(137,128){1}
//: {2}(139,126)(183,126){3}
//: {4}(137,124)(137,87)(95,87){5}
output c;    //: /sn:0 /dp:1 {0}(204,164)(243,164){1}
//: enddecls

  //: output g4 (s) @(238,129) /sn:0 /w:[ 1 ]
  //: input g3 (b) @(92,103) /sn:0 /w:[ 0 ]
  //: input g2 (a) @(93,87) /sn:0 /w:[ 5 ]
  and g1 (.I0(a), .I1(b), .Z(c));   //: @(194,164) /sn:0 /delay:" 5" /w:[ 0 5 0 ]
  //: joint g6 (b) @(125, 131) /w:[ 2 1 -1 4 ]
  //: joint g7 (a) @(137, 126) /w:[ 2 4 -1 1 ]
  //: output g5 (c) @(240,164) /sn:0 /w:[ 1 ]
  xor g0 (.I0(a), .I1(b), .Z(s));   //: @(194,129) /sn:0 /delay:" 6" /w:[ 3 3 0 ]

endmodule

module FA(c_out, s, c_in, b, a);
//: interface  /sz:(57, 40) /bd:[ Ti0>a(41/57) Ti1>b(21/57) Ri0>c_in(19/40) Lo0<c_out(19/40) Bo0<s(29/57) ]
input b;    //: /sn:0 /dp:1 {0}(240,94)(203,94)(203,34){1}
output c_out;    //: /sn:0 /dp:1 {0}(404,147)(427,147){1}
input c_in;    //: /sn:0 {0}(299,37)(299,84)(333,84){1}
output s;    //: /sn:0 {0}(429,93)(379,93){1}
input a;    //: /sn:0 {0}(187,34)(187,113)(240,113){1}
wire w4;    //: /sn:0 /dp:1 {0}(383,149)(261,149)(261,126){1}
wire w0;    //: /sn:0 /dp:1 {0}(383,144)(354,144)(354,116){1}
wire w5;    //: /sn:0 {0}(286,103)(333,103){1}
//: enddecls

  //: output g4 (c_out) @(424,147) /sn:0 /w:[ 1 ]
  //: output g3 (s) @(426,93) /sn:0 /w:[ 0 ]
  //: input g2 (c_in) @(299,35) /sn:0 /R:3 /w:[ 0 ]
  //: input g1 (b) @(203,32) /sn:0 /R:3 /w:[ 1 ]
  or g7 (.I0(w0), .I1(w4), .Z(c_out));   //: @(394,147) /sn:0 /delay:" 5" /w:[ 0 0 0 ]
  HA g14 (.b(b), .a(a), .c(w4), .s(w5));   //: @(241, 81) /sz:(44, 44) /sn:0 /p:[ Li0>0 Li1>1 Bo0<1 Ro0<0 ]
  HA g15 (.b(c_in), .a(w5), .c(w0), .s(s));   //: @(334, 71) /sz:(44, 44) /sn:0 /p:[ Li0>1 Li1>1 Bo0<1 Ro0<1 ]
  //: input g0 (a) @(187,32) /sn:0 /R:3 /w:[ 0 ]

endmodule

module main;    //: root_module
wire [3:0] w0;    //: /sn:0 /dp:1 {0}(431,185)(431,124)(382,124)(382,76){1}
wire [7:0] w3;    //: /sn:0 {0}(325,294)(325,346)(447,346)(447,260){1}
wire [3:0] w2;    //: /sn:0 {0}(511,76)(511,123)(466,123)(466,185){1}
//: enddecls

  //: dip g3 (w2) @(511,66) /sn:0 /w:[ 0 ] /st:15
  //: dip g2 (w0) @(382,66) /sn:0 /w:[ 1 ] /st:15
  led g1 (.I(w3));   //: @(325,287) /sn:0 /w:[ 0 ] /type:3
  RCA4bits g0 (.b(w2), .a(w0), .s(w3));   //: @(409, 186) /sz:(77, 73) /sn:0 /p:[ Ti0>1 Ti1>0 Bo0<1 ]

endmodule
